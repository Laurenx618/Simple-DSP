`timescale 1ns/1ps
`default_nettype none
`include "hdl/register.sv"

//////////////////////////////////////////////////////////////////////////////////////
// This is the main Verilog hdl file automatically generated from filter.py
// The block diagram of the FIR filter we build can be accessed in this github repo
//////////////////////////////////////////////////////////////////////////////////////

module fir(clk, rst, ena, filter_select, sample, out);

    input wire clk, rst, ena;
    input wire filter_select;
    input wire [15:0] sample;
    output logic [32:0] out;


    ////// TAP COEFFICIENTS //////
    logic signed [15:0] tap0, tap1, tap2, tap3, tap4, tap5, tap6, tap7, tap8, tap9, tap10, tap11, tap12, tap13, tap14, tap15, tap16, tap17, tap18, tap19, tap20, tap21, tap22, tap23, tap24, tap25, tap26, tap27, tap28, tap29, tap30, tap31, tap32, tap33, tap34, tap35, tap36, tap37, tap38, tap39, tap40, tap41, tap42, tap43, tap44, tap45, tap46, tap47, tap48, tap49, tap50, tap51, tap52, tap53, tap54, tap55, tap56, tap57, tap58, tap59, tap60, tap61, tap62, tap63, tap64, tap65, tap66, tap67, tap68, tap69, tap70, tap71, tap72, tap73, tap74;
    mux2_16 tap0_mux (.a({-16'sd42, 16'sd42}), .s(filter_select), .y(tap0);
    mux2_16 tap1_mux (.a({-16'sd27, 16'sd27}), .s(filter_select), .y(tap1);
    mux2_16 tap2_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap2);
    mux2_16 tap3_mux (.a({16'sd34, -16'sd34}), .s(filter_select), .y(tap3);
    mux2_16 tap4_mux (.a({16'sd63, -16'sd63}), .s(filter_select), .y(tap4);
    mux2_16 tap5_mux (.a({16'sd74, -16'sd74}), .s(filter_select), .y(tap5);
    mux2_16 tap6_mux (.a({16'sd54, -16'sd54}), .s(filter_select), .y(tap6);
    mux2_16 tap7_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap7);
    mux2_16 tap8_mux (.a({-16'sd76, 16'sd77}), .s(filter_select), .y(tap8);
    mux2_16 tap9_mux (.a({-16'sd147, 16'sd147}), .s(filter_select), .y(tap9);
    mux2_16 tap10_mux (.a({-16'sd173, 16'sd173}), .s(filter_select), .y(tap10);
    mux2_16 tap11_mux (.a({-16'sd125, 16'sd125}), .s(filter_select), .y(tap11);
    mux2_16 tap12_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap12);
    mux2_16 tap13_mux (.a({16'sd170, -16'sd170}), .s(filter_select), .y(tap13);
    mux2_16 tap14_mux (.a({16'sd317, -16'sd318}), .s(filter_select), .y(tap14);
    mux2_16 tap15_mux (.a({16'sd365, -16'sd365}), .s(filter_select), .y(tap15);
    mux2_16 tap16_mux (.a({16'sd258, -16'sd258}), .s(filter_select), .y(tap16);
    mux2_16 tap17_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap17);
    mux2_16 tap18_mux (.a({-16'sd335, 16'sd336}), .s(filter_select), .y(tap18);
    mux2_16 tap19_mux (.a({-16'sd616, 16'sd617}), .s(filter_select), .y(tap19);
    mux2_16 tap20_mux (.a({-16'sd698, 16'sd698}), .s(filter_select), .y(tap20);
    mux2_16 tap21_mux (.a({-16'sd488, 16'sd488}), .s(filter_select), .y(tap21);
    mux2_16 tap22_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap22);
    mux2_16 tap23_mux (.a({16'sd623, -16'sd623}), .s(filter_select), .y(tap23);
    mux2_16 tap24_mux (.a({16'sd1140, -16'sd1140}), .s(filter_select), .y(tap24);
    mux2_16 tap25_mux (.a({16'sd1291, -16'sd1292}), .s(filter_select), .y(tap25);
    mux2_16 tap26_mux (.a({16'sd906, -16'sd907}), .s(filter_select), .y(tap26);
    mux2_16 tap27_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap27);
    mux2_16 tap28_mux (.a({-16'sd1188, 16'sd1189}), .s(filter_select), .y(tap28);
    mux2_16 tap29_mux (.a({-16'sd2226, 16'sd2228}), .s(filter_select), .y(tap29);
    mux2_16 tap30_mux (.a({-16'sd2610, 16'sd2612}), .s(filter_select), .y(tap30);
    mux2_16 tap31_mux (.a({-16'sd1924, 16'sd1925}), .s(filter_select), .y(tap31);
    mux2_16 tap32_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap32);
    mux2_16 tap33_mux (.a({16'sd2984, -16'sd2986}), .s(filter_select), .y(tap33);
    mux2_16 tap34_mux (.a({16'sd6515, -16'sd6519}), .s(filter_select), .y(tap34);
    mux2_16 tap35_mux (.a({16'sd9854, -16'sd9861}), .s(filter_select), .y(tap35);
    mux2_16 tap36_mux (.a({16'sd12241, -16'sd12250}), .s(filter_select), .y(tap36);
    mux2_16 tap37_mux (.a({16'sd13107, 16'sd52466}), .s(filter_select), .y(tap37);
    mux2_16 tap38_mux (.a({16'sd12241, -16'sd12250}), .s(filter_select), .y(tap38);
    mux2_16 tap39_mux (.a({16'sd9854, -16'sd9861}), .s(filter_select), .y(tap39);
    mux2_16 tap40_mux (.a({16'sd6515, -16'sd6519}), .s(filter_select), .y(tap40);
    mux2_16 tap41_mux (.a({16'sd2984, -16'sd2986}), .s(filter_select), .y(tap41);
    mux2_16 tap42_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap42);
    mux2_16 tap43_mux (.a({-16'sd1924, 16'sd1925}), .s(filter_select), .y(tap43);
    mux2_16 tap44_mux (.a({-16'sd2610, 16'sd2612}), .s(filter_select), .y(tap44);
    mux2_16 tap45_mux (.a({-16'sd2226, 16'sd2228}), .s(filter_select), .y(tap45);
    mux2_16 tap46_mux (.a({-16'sd1188, 16'sd1189}), .s(filter_select), .y(tap46);
    mux2_16 tap47_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap47);
    mux2_16 tap48_mux (.a({16'sd906, -16'sd907}), .s(filter_select), .y(tap48);
    mux2_16 tap49_mux (.a({16'sd1291, -16'sd1292}), .s(filter_select), .y(tap49);
    mux2_16 tap50_mux (.a({16'sd1140, -16'sd1140}), .s(filter_select), .y(tap50);
    mux2_16 tap51_mux (.a({16'sd623, -16'sd623}), .s(filter_select), .y(tap51);
    mux2_16 tap52_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap52);
    mux2_16 tap53_mux (.a({-16'sd488, 16'sd488}), .s(filter_select), .y(tap53);
    mux2_16 tap54_mux (.a({-16'sd698, 16'sd698}), .s(filter_select), .y(tap54);
    mux2_16 tap55_mux (.a({-16'sd616, 16'sd617}), .s(filter_select), .y(tap55);
    mux2_16 tap56_mux (.a({-16'sd335, 16'sd336}), .s(filter_select), .y(tap56);
    mux2_16 tap57_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap57);
    mux2_16 tap58_mux (.a({16'sd258, -16'sd258}), .s(filter_select), .y(tap58);
    mux2_16 tap59_mux (.a({16'sd365, -16'sd365}), .s(filter_select), .y(tap59);
    mux2_16 tap60_mux (.a({16'sd317, -16'sd318}), .s(filter_select), .y(tap60);
    mux2_16 tap61_mux (.a({16'sd170, -16'sd170}), .s(filter_select), .y(tap61);
    mux2_16 tap62_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap62);
    mux2_16 tap63_mux (.a({-16'sd125, 16'sd125}), .s(filter_select), .y(tap63);
    mux2_16 tap64_mux (.a({-16'sd173, 16'sd173}), .s(filter_select), .y(tap64);
    mux2_16 tap65_mux (.a({-16'sd147, 16'sd147}), .s(filter_select), .y(tap65);
    mux2_16 tap66_mux (.a({-16'sd76, 16'sd77}), .s(filter_select), .y(tap66);
    mux2_16 tap67_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap67);
    mux2_16 tap68_mux (.a({16'sd54, -16'sd54}), .s(filter_select), .y(tap68);
    mux2_16 tap69_mux (.a({16'sd74, -16'sd74}), .s(filter_select), .y(tap69);
    mux2_16 tap70_mux (.a({16'sd63, -16'sd63}), .s(filter_select), .y(tap70);
    mux2_16 tap71_mux (.a({16'sd34, -16'sd34}), .s(filter_select), .y(tap71);
    mux2_16 tap72_mux (.a({16'sd0, 16'sd0}), .s(filter_select), .y(tap72);
    mux2_16 tap73_mux (.a({-16'sd27, 16'sd27}), .s(filter_select), .y(tap73);
    mux2_16 tap74_mux (.a({-16'sd42, 16'sd42}), .s(filter_select), .y(tap74);


    ////// SAMPLE SHIFT REGISTER //////
    logic signed [15:0] buf0, buf1, buf2, buf3, buf4, buf5, buf6, buf7, buf8, buf9, buf10, buf11, buf12, buf13, buf14, buf15, buf16, buf17, buf18, buf19, buf20, buf21, buf22, buf23, buf24, buf25, buf26, buf27, buf28, buf29, buf30, buf31, buf32, buf33, buf34, buf35, buf36, buf37, buf38, buf39, buf40, buf41, buf42, buf43, buf44, buf45, buf46, buf47, buf48, buf49, buf50, buf51, buf52, buf53, buf54, buf55, buf56, buf57, buf58, buf59, buf60, buf61, buf62, buf63, buf64, buf65, buf66, buf67, buf68, buf69, buf70, buf71, buf72, buf73, buf74;
    register #(.N(16)) buffer0(.clk(clk), .ena(ena), .rst(rst), .d(sample), .q(buf0));
    register #(.N(16)) buffer1(.clk(clk), .ena(ena), .rst(rst), .d(buf0), .q(buf1));
    register #(.N(16)) buffer2(.clk(clk), .ena(ena), .rst(rst), .d(buf1), .q(buf2));
    register #(.N(16)) buffer3(.clk(clk), .ena(ena), .rst(rst), .d(buf2), .q(buf3));
    register #(.N(16)) buffer4(.clk(clk), .ena(ena), .rst(rst), .d(buf3), .q(buf4));
    register #(.N(16)) buffer5(.clk(clk), .ena(ena), .rst(rst), .d(buf4), .q(buf5));
    register #(.N(16)) buffer6(.clk(clk), .ena(ena), .rst(rst), .d(buf5), .q(buf6));
    register #(.N(16)) buffer7(.clk(clk), .ena(ena), .rst(rst), .d(buf6), .q(buf7));
    register #(.N(16)) buffer8(.clk(clk), .ena(ena), .rst(rst), .d(buf7), .q(buf8));
    register #(.N(16)) buffer9(.clk(clk), .ena(ena), .rst(rst), .d(buf8), .q(buf9));
    register #(.N(16)) buffer10(.clk(clk), .ena(ena), .rst(rst), .d(buf9), .q(buf10));
    register #(.N(16)) buffer11(.clk(clk), .ena(ena), .rst(rst), .d(buf10), .q(buf11));
    register #(.N(16)) buffer12(.clk(clk), .ena(ena), .rst(rst), .d(buf11), .q(buf12));
    register #(.N(16)) buffer13(.clk(clk), .ena(ena), .rst(rst), .d(buf12), .q(buf13));
    register #(.N(16)) buffer14(.clk(clk), .ena(ena), .rst(rst), .d(buf13), .q(buf14));
    register #(.N(16)) buffer15(.clk(clk), .ena(ena), .rst(rst), .d(buf14), .q(buf15));
    register #(.N(16)) buffer16(.clk(clk), .ena(ena), .rst(rst), .d(buf15), .q(buf16));
    register #(.N(16)) buffer17(.clk(clk), .ena(ena), .rst(rst), .d(buf16), .q(buf17));
    register #(.N(16)) buffer18(.clk(clk), .ena(ena), .rst(rst), .d(buf17), .q(buf18));
    register #(.N(16)) buffer19(.clk(clk), .ena(ena), .rst(rst), .d(buf18), .q(buf19));
    register #(.N(16)) buffer20(.clk(clk), .ena(ena), .rst(rst), .d(buf19), .q(buf20));
    register #(.N(16)) buffer21(.clk(clk), .ena(ena), .rst(rst), .d(buf20), .q(buf21));
    register #(.N(16)) buffer22(.clk(clk), .ena(ena), .rst(rst), .d(buf21), .q(buf22));
    register #(.N(16)) buffer23(.clk(clk), .ena(ena), .rst(rst), .d(buf22), .q(buf23));
    register #(.N(16)) buffer24(.clk(clk), .ena(ena), .rst(rst), .d(buf23), .q(buf24));
    register #(.N(16)) buffer25(.clk(clk), .ena(ena), .rst(rst), .d(buf24), .q(buf25));
    register #(.N(16)) buffer26(.clk(clk), .ena(ena), .rst(rst), .d(buf25), .q(buf26));
    register #(.N(16)) buffer27(.clk(clk), .ena(ena), .rst(rst), .d(buf26), .q(buf27));
    register #(.N(16)) buffer28(.clk(clk), .ena(ena), .rst(rst), .d(buf27), .q(buf28));
    register #(.N(16)) buffer29(.clk(clk), .ena(ena), .rst(rst), .d(buf28), .q(buf29));
    register #(.N(16)) buffer30(.clk(clk), .ena(ena), .rst(rst), .d(buf29), .q(buf30));
    register #(.N(16)) buffer31(.clk(clk), .ena(ena), .rst(rst), .d(buf30), .q(buf31));
    register #(.N(16)) buffer32(.clk(clk), .ena(ena), .rst(rst), .d(buf31), .q(buf32));
    register #(.N(16)) buffer33(.clk(clk), .ena(ena), .rst(rst), .d(buf32), .q(buf33));
    register #(.N(16)) buffer34(.clk(clk), .ena(ena), .rst(rst), .d(buf33), .q(buf34));
    register #(.N(16)) buffer35(.clk(clk), .ena(ena), .rst(rst), .d(buf34), .q(buf35));
    register #(.N(16)) buffer36(.clk(clk), .ena(ena), .rst(rst), .d(buf35), .q(buf36));
    register #(.N(16)) buffer37(.clk(clk), .ena(ena), .rst(rst), .d(buf36), .q(buf37));
    register #(.N(16)) buffer38(.clk(clk), .ena(ena), .rst(rst), .d(buf37), .q(buf38));
    register #(.N(16)) buffer39(.clk(clk), .ena(ena), .rst(rst), .d(buf38), .q(buf39));
    register #(.N(16)) buffer40(.clk(clk), .ena(ena), .rst(rst), .d(buf39), .q(buf40));
    register #(.N(16)) buffer41(.clk(clk), .ena(ena), .rst(rst), .d(buf40), .q(buf41));
    register #(.N(16)) buffer42(.clk(clk), .ena(ena), .rst(rst), .d(buf41), .q(buf42));
    register #(.N(16)) buffer43(.clk(clk), .ena(ena), .rst(rst), .d(buf42), .q(buf43));
    register #(.N(16)) buffer44(.clk(clk), .ena(ena), .rst(rst), .d(buf43), .q(buf44));
    register #(.N(16)) buffer45(.clk(clk), .ena(ena), .rst(rst), .d(buf44), .q(buf45));
    register #(.N(16)) buffer46(.clk(clk), .ena(ena), .rst(rst), .d(buf45), .q(buf46));
    register #(.N(16)) buffer47(.clk(clk), .ena(ena), .rst(rst), .d(buf46), .q(buf47));
    register #(.N(16)) buffer48(.clk(clk), .ena(ena), .rst(rst), .d(buf47), .q(buf48));
    register #(.N(16)) buffer49(.clk(clk), .ena(ena), .rst(rst), .d(buf48), .q(buf49));
    register #(.N(16)) buffer50(.clk(clk), .ena(ena), .rst(rst), .d(buf49), .q(buf50));
    register #(.N(16)) buffer51(.clk(clk), .ena(ena), .rst(rst), .d(buf50), .q(buf51));
    register #(.N(16)) buffer52(.clk(clk), .ena(ena), .rst(rst), .d(buf51), .q(buf52));
    register #(.N(16)) buffer53(.clk(clk), .ena(ena), .rst(rst), .d(buf52), .q(buf53));
    register #(.N(16)) buffer54(.clk(clk), .ena(ena), .rst(rst), .d(buf53), .q(buf54));
    register #(.N(16)) buffer55(.clk(clk), .ena(ena), .rst(rst), .d(buf54), .q(buf55));
    register #(.N(16)) buffer56(.clk(clk), .ena(ena), .rst(rst), .d(buf55), .q(buf56));
    register #(.N(16)) buffer57(.clk(clk), .ena(ena), .rst(rst), .d(buf56), .q(buf57));
    register #(.N(16)) buffer58(.clk(clk), .ena(ena), .rst(rst), .d(buf57), .q(buf58));
    register #(.N(16)) buffer59(.clk(clk), .ena(ena), .rst(rst), .d(buf58), .q(buf59));
    register #(.N(16)) buffer60(.clk(clk), .ena(ena), .rst(rst), .d(buf59), .q(buf60));
    register #(.N(16)) buffer61(.clk(clk), .ena(ena), .rst(rst), .d(buf60), .q(buf61));
    register #(.N(16)) buffer62(.clk(clk), .ena(ena), .rst(rst), .d(buf61), .q(buf62));
    register #(.N(16)) buffer63(.clk(clk), .ena(ena), .rst(rst), .d(buf62), .q(buf63));
    register #(.N(16)) buffer64(.clk(clk), .ena(ena), .rst(rst), .d(buf63), .q(buf64));
    register #(.N(16)) buffer65(.clk(clk), .ena(ena), .rst(rst), .d(buf64), .q(buf65));
    register #(.N(16)) buffer66(.clk(clk), .ena(ena), .rst(rst), .d(buf65), .q(buf66));
    register #(.N(16)) buffer67(.clk(clk), .ena(ena), .rst(rst), .d(buf66), .q(buf67));
    register #(.N(16)) buffer68(.clk(clk), .ena(ena), .rst(rst), .d(buf67), .q(buf68));
    register #(.N(16)) buffer69(.clk(clk), .ena(ena), .rst(rst), .d(buf68), .q(buf69));
    register #(.N(16)) buffer70(.clk(clk), .ena(ena), .rst(rst), .d(buf69), .q(buf70));
    register #(.N(16)) buffer71(.clk(clk), .ena(ena), .rst(rst), .d(buf70), .q(buf71));
    register #(.N(16)) buffer72(.clk(clk), .ena(ena), .rst(rst), .d(buf71), .q(buf72));
    register #(.N(16)) buffer73(.clk(clk), .ena(ena), .rst(rst), .d(buf72), .q(buf73));
    register #(.N(16)) buffer74(.clk(clk), .ena(ena), .rst(rst), .d(buf73), .q(buf74));


    ////// LINEAR COMBINATION SAMPLES WITH TAPS //////
    logic signed [31:0] multiplied0, multiplied1, multiplied2, multiplied3, multiplied4, multiplied5, multiplied6, multiplied7, multiplied8, multiplied9, multiplied10, multiplied11, multiplied12, multiplied13, multiplied14, multiplied15, multiplied16, multiplied17, multiplied18, multiplied19, multiplied20, multiplied21, multiplied22, multiplied23, multiplied24, multiplied25, multiplied26, multiplied27, multiplied28, multiplied29, multiplied30, multiplied31, multiplied32, multiplied33, multiplied34, multiplied35, multiplied36, multiplied37, multiplied38, multiplied39, multiplied40, multiplied41, multiplied42, multiplied43, multiplied44, multiplied45, multiplied46, multiplied47, multiplied48, multiplied49, multiplied50, multiplied51, multiplied52, multiplied53, multiplied54, multiplied55, multiplied56, multiplied57, multiplied58, multiplied59, multiplied60, multiplied61, multiplied62, multiplied63, multiplied64, multiplied65, multiplied66, multiplied67, multiplied68, multiplied69, multiplied70, multiplied71, multiplied72, multiplied73, multiplied74;
    always_comb multiplied0 = buf0 * tap0;
    always_comb multiplied1 = buf1 * tap1;
    always_comb multiplied2 = buf2 * tap2;
    always_comb multiplied3 = buf3 * tap3;
    always_comb multiplied4 = buf4 * tap4;
    always_comb multiplied5 = buf5 * tap5;
    always_comb multiplied6 = buf6 * tap6;
    always_comb multiplied7 = buf7 * tap7;
    always_comb multiplied8 = buf8 * tap8;
    always_comb multiplied9 = buf9 * tap9;
    always_comb multiplied10 = buf10 * tap10;
    always_comb multiplied11 = buf11 * tap11;
    always_comb multiplied12 = buf12 * tap12;
    always_comb multiplied13 = buf13 * tap13;
    always_comb multiplied14 = buf14 * tap14;
    always_comb multiplied15 = buf15 * tap15;
    always_comb multiplied16 = buf16 * tap16;
    always_comb multiplied17 = buf17 * tap17;
    always_comb multiplied18 = buf18 * tap18;
    always_comb multiplied19 = buf19 * tap19;
    always_comb multiplied20 = buf20 * tap20;
    always_comb multiplied21 = buf21 * tap21;
    always_comb multiplied22 = buf22 * tap22;
    always_comb multiplied23 = buf23 * tap23;
    always_comb multiplied24 = buf24 * tap24;
    always_comb multiplied25 = buf25 * tap25;
    always_comb multiplied26 = buf26 * tap26;
    always_comb multiplied27 = buf27 * tap27;
    always_comb multiplied28 = buf28 * tap28;
    always_comb multiplied29 = buf29 * tap29;
    always_comb multiplied30 = buf30 * tap30;
    always_comb multiplied31 = buf31 * tap31;
    always_comb multiplied32 = buf32 * tap32;
    always_comb multiplied33 = buf33 * tap33;
    always_comb multiplied34 = buf34 * tap34;
    always_comb multiplied35 = buf35 * tap35;
    always_comb multiplied36 = buf36 * tap36;
    always_comb multiplied37 = buf37 * tap37;
    always_comb multiplied38 = buf38 * tap38;
    always_comb multiplied39 = buf39 * tap39;
    always_comb multiplied40 = buf40 * tap40;
    always_comb multiplied41 = buf41 * tap41;
    always_comb multiplied42 = buf42 * tap42;
    always_comb multiplied43 = buf43 * tap43;
    always_comb multiplied44 = buf44 * tap44;
    always_comb multiplied45 = buf45 * tap45;
    always_comb multiplied46 = buf46 * tap46;
    always_comb multiplied47 = buf47 * tap47;
    always_comb multiplied48 = buf48 * tap48;
    always_comb multiplied49 = buf49 * tap49;
    always_comb multiplied50 = buf50 * tap50;
    always_comb multiplied51 = buf51 * tap51;
    always_comb multiplied52 = buf52 * tap52;
    always_comb multiplied53 = buf53 * tap53;
    always_comb multiplied54 = buf54 * tap54;
    always_comb multiplied55 = buf55 * tap55;
    always_comb multiplied56 = buf56 * tap56;
    always_comb multiplied57 = buf57 * tap57;
    always_comb multiplied58 = buf58 * tap58;
    always_comb multiplied59 = buf59 * tap59;
    always_comb multiplied60 = buf60 * tap60;
    always_comb multiplied61 = buf61 * tap61;
    always_comb multiplied62 = buf62 * tap62;
    always_comb multiplied63 = buf63 * tap63;
    always_comb multiplied64 = buf64 * tap64;
    always_comb multiplied65 = buf65 * tap65;
    always_comb multiplied66 = buf66 * tap66;
    always_comb multiplied67 = buf67 * tap67;
    always_comb multiplied68 = buf68 * tap68;
    always_comb multiplied69 = buf69 * tap69;
    always_comb multiplied70 = buf70 * tap70;
    always_comb multiplied71 = buf71 * tap71;
    always_comb multiplied72 = buf72 * tap72;
    always_comb multiplied73 = buf73 * tap73;
    always_comb multiplied74 = buf74 * tap74;

    always_comb out = multiplied0 + multiplied1 + multiplied2 + multiplied3 + multiplied4 + multiplied5 + multiplied6 + multiplied7 + multiplied8 + multiplied9 + multiplied10 + multiplied11 + multiplied12 + multiplied13 + multiplied14 + multiplied15 + multiplied16 + multiplied17 + multiplied18 + multiplied19 + multiplied20 + multiplied21 + multiplied22 + multiplied23 + multiplied24 + multiplied25 + multiplied26 + multiplied27 + multiplied28 + multiplied29 + multiplied30 + multiplied31 + multiplied32 + multiplied33 + multiplied34 + multiplied35 + multiplied36 + multiplied37 + multiplied38 + multiplied39 + multiplied40 + multiplied41 + multiplied42 + multiplied43 + multiplied44 + multiplied45 + multiplied46 + multiplied47 + multiplied48 + multiplied49 + multiplied50 + multiplied51 + multiplied52 + multiplied53 + multiplied54 + multiplied55 + multiplied56 + multiplied57 + multiplied58 + multiplied59 + multiplied60 + multiplied61 + multiplied62 + multiplied63 + multiplied64 + multiplied65 + multiplied66 + multiplied67 + multiplied68 + multiplied69 + multiplied70 + multiplied71 + multiplied72 + multiplied73 + multiplied74;

endmodule