`timescale 1ns/1ps
`default_nettype none

module test_fir;
int errors = 0;

logic rst;
logic clk;
logic shift_ena;
logic [15:0] next_sample;
logic [38:0] out;

logic [8:0] counter;
logic [38:0] correct_out;

// integer samples [399:0];
// time correct_outputs [399:0];

integer test[7:0] = '{26, 40, 32, 18, 50, 0, 20, 12};


// integer xyzzy[7:0] = '{26, 40, 32, 18, 50, 0, 20, 12};

logic [15:0] samples [399:0] = '{72200, 90564, 84560, 69249, 61880, 62782, 68570, 81332, 94609, 90928, 68018, 50830, 60149, 82167, 87989, 73243, 57675, 52510, 51258, 50538, 55715, 62361, 55290, 34526, 21916, 30203, 43308, 41391, 29511, 24186, 25102, 21159, 15385, 20309, 32017, 32431, 19016, 10144, 15839, 24055, 24052, 23069, 27703, 27689, 15133, 4539, 13068, 30953, 33500, 17189, 2083, 285, 3981, 6034, 9679, 11979, 273, -23603, -35588, -21648, -2036, -5176, -29137, -48491, -50637, -44308, -37770, -31734, -32851, -49977, -72284, -73939, -50365, -30053, -37381, -60647, -72199, -65414, -53639, -44751, -38284, -39913, -54997, -69881, -63259, -39071, -26151, -38780, -58084, -61974, -53912, -48621, -47214, -44413, -46378, -60060, -73625, -69785, -54562, -50811, -63842, -75484, -74877, -72574, -76889, -78285, -69917, -64582, -74259, -87402, -85623, -72412, -65348, -67389, -67272, -63934, -67143, -73576, -66462, -45189, -32841, -43136, -58894, -57455, -41512, -28654, -24131, -22699, -26315, -37964, -44563, -30123, -5142, 803, -19940, -41141, -39240, -21920, -9767, -8381, -12995, -23823, -38106, -39920, -19831, 2908, 475, -24053, -39415, -28863, -8252, 2297, 2573, -201, -6524, -13625, -7621, 15524, 34841, 29802, 11438, 7624, 23788, 40026, 44162, 44243, 46388, 44119, 37264, 39659, 55722, 67626, 60806, 47107, 45709, 53871, 56109, 52444, 54953, 61471, 57052, 42284, 36632, 47857, 59327, 56694, 47929, 45194, 44894, 41038, 42346, 56495, 69175, 61417, 41542, 36777, 54359, 73163, 76108, 69276, 63563, 59005, 56979, 67306, 88359, 97492, 80076, 55594, 54275, 75927, 93004, 89641, 75718, 63820, 55526, 53710, 64926, 80774, 78167, 51607, 27679, 31352, 51987, 60659, 49618, 34417, 25441, 20213, 20188, 30859, 43109, 37752, 15623, 2352, 13036, 30861, 33647, 24387, 19070, 19062, 16004, 13667, 21902, 33662, 31294, 15725, 7297, 14211, 21534, 18099, 13075, 14897, 13663, 496, -11880, -7586, 4738, 3732, -12195, -25387, -28104, -29130, -31812, -28790, -22976, -30556, -52992, -66681, -55179, -35119, -33006, -49211, -63552, -66259, -62817, -55393, -42605, -35234, -47762, -70903, -75619, -52851, -28929, -29994, -49024, -62122, -61365, -54274, -44363, -33227, -32705, -51548, -73528, -72226, -48969, -34001, -45172, -66553, -75999, -73381, -69255, -64503, -58211, -60628, -77811, -93445, -87555, -67699, -59904, -70989, -82065, -80488, -75171, -74270, -70330, -59084, -53206, -61601, -70581, -63552, -47489, -40689, -43481, -42192, -36149, -37264, -43871, -39331, -21535, -11103, -20502, -34650, -34814, -24749, -18246, -15960, -12598, -14486, -28329, -40490, -31319, -7952, 657, -15831, -35487, -36772, -24243, -12673, -5511, -2311, -9437, -25482, -30192, -9126, 19530, 24844, 5447, -9852, -2557, 16510, 30895, 38336, 39908, 31520, 18804, 21432, 45866, 68469, 64470, 42914, 32951, 43357, 57234, 62299, 62881, 61428, 52203, 39608, 40547, 57687, 69331, 59531, 42018, 38357, 46595, 50475, 48395, 50949, 56230, 51666, 39761, 38568, 52410, 63591, 60569, 54303, 56340, 59885, 56962, 57159};
logic [38:0] correct_outputs [399:0] = '{-680344, -1249027, -729189, 1604747, 5510102, 9517597, 11225695, 8257649, -193474, -12036352, -22348746, -25225238, -16561402, 3491148, 29339678, 50756621, 56169119, 37863337, -3036453, -54530355, -96273242, -106458679, -71194131, 6905391, 105038314, 184675544, 204221742, 136129330, -17532302, -217019524, -388544939, -440467321, -288384022, 118584483, 779191628, 1635563348, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2119050508, 1961578198, 1825613808, 1711726412, 1618520094, 1543913620, 1486144420, 1443869537, 1415644487, 1399583439, 1393463392, 1395334482, 1401729440, 1409349257, 1415045527, 1415850343, 1408712506, 1390536666, 1358577801, 1310619698, 1244769489, 1159378250, 1053322259, 926173231, 777959263, 608969735, 420003136, 212650657, -10913061, -248349975, -497174709, -754468102, -1016886292, -1281003119, -1543457205, -1800804872, -2049565754, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116424109, -1966200130, -1833456980, -1719204103, -1623656724, -1546414429, -1486748438, -1443526511, -1415026426, -1399085387, -1393370079, -1395295928, -1401790068, -1409464270, -1415100177, -1415786123, -1408603216, -1390497512, -1358629108, -1310688480, -1244798133, -1159370150, -1053293395, -926128433, -777925344, -608988455, -420066199, -212691504, 10934638, 248397668, 497197646, 754467482, 1016883018, 1280984437, 1543410748, 1800774184, 2049604907, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2116432099, 1966254228, 1833495929, 1719199916, 1623634864, 1546392840, 1486718012, 1443502820, 1415054996, 1399162709, 1393414651, 1395245950, 1401693470, 1409422554, 1415147310, 1415868176, 1408654856, 1390489290, 1358560455, 1310596159, 1244764317, 1159451978, 1053428891, 926175129, 777824466, 608843488, 420023277, 212780111, -10808148, -248337736, -497242634, -754585812, -1016987672, -1280976052, -1543274751, -1800632613, -2049607436, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116288505, -1966208814, -1833573049, -1719323701, -1623710967, -1546362187, -1486591395, -1443380596, -1415061729, -1399309517, -1393558099, -1395236836, -1401547290, -1409293513, -1415149926, -1415976828, -1408766703, -1390523934, -1358496187, -1310475479, -1244686307, -1159499955, -1053567883, -926264615, -777772732, -608714815, -419953035, -212818149, 10723054, 248279976, 497238088, 754630761, 1017059437, 1281019096, 1543239093, 1800546637, 2049562238};
// always_comb samples = '{72200, 90564, 84560, 69249, 61880, 62782, 68570, 81332, 94609, 90928, 68018, 50830, 60149, 82167, 87989, 73243, 57675, 52510, 51258, 50538, 55715, 62361, 55290, 34526, 21916, 30203, 43308, 41391, 29511, 24186, 25102, 21159, 15385, 20309, 32017, 32431, 19016, 10144, 15839, 24055, 24052, 23069, 27703, 27689, 15133, 4539, 13068, 30953, 33500, 17189, 2083, 285, 3981, 6034, 9679, 11979, 273, -23603, -35588, -21648, -2036, -5176, -29137, -48491, -50637, -44308, -37770, -31734, -32851, -49977, -72284, -73939, -50365, -30053, -37381, -60647, -72199, -65414, -53639, -44751, -38284, -39913, -54997, -69881, -63259, -39071, -26151, -38780, -58084, -61974, -53912, -48621, -47214, -44413, -46378, -60060, -73625, -69785, -54562, -50811, -63842, -75484, -74877, -72574, -76889, -78285, -69917, -64582, -74259, -87402, -85623, -72412, -65348, -67389, -67272, -63934, -67143, -73576, -66462, -45189, -32841, -43136, -58894, -57455, -41512, -28654, -24131, -22699, -26315, -37964, -44563, -30123, -5142, 803, -19940, -41141, -39240, -21920, -9767, -8381, -12995, -23823, -38106, -39920, -19831, 2908, 475, -24053, -39415, -28863, -8252, 2297, 2573, -201, -6524, -13625, -7621, 15524, 34841, 29802, 11438, 7624, 23788, 40026, 44162, 44243, 46388, 44119, 37264, 39659, 55722, 67626, 60806, 47107, 45709, 53871, 56109, 52444, 54953, 61471, 57052, 42284, 36632, 47857, 59327, 56694, 47929, 45194, 44894, 41038, 42346, 56495, 69175, 61417, 41542, 36777, 54359, 73163, 76108, 69276, 63563, 59005, 56979, 67306, 88359, 97492, 80076, 55594, 54275, 75927, 93004, 89641, 75718, 63820, 55526, 53710, 64926, 80774, 78167, 51607, 27679, 31352, 51987, 60659, 49618, 34417, 25441, 20213, 20188, 30859, 43109, 37752, 15623, 2352, 13036, 30861, 33647, 24387, 19070, 19062, 16004, 13667, 21902, 33662, 31294, 15725, 7297, 14211, 21534, 18099, 13075, 14897, 13663, 496, -11880, -7586, 4738, 3732, -12195, -25387, -28104, -29130, -31812, -28790, -22976, -30556, -52992, -66681, -55179, -35119, -33006, -49211, -63552, -66259, -62817, -55393, -42605, -35234, -47762, -70903, -75619, -52851, -28929, -29994, -49024, -62122, -61365, -54274, -44363, -33227, -32705, -51548, -73528, -72226, -48969, -34001, -45172, -66553, -75999, -73381, -69255, -64503, -58211, -60628, -77811, -93445, -87555, -67699, -59904, -70989, -82065, -80488, -75171, -74270, -70330, -59084, -53206, -61601, -70581, -63552, -47489, -40689, -43481, -42192, -36149, -37264, -43871, -39331, -21535, -11103, -20502, -34650, -34814, -24749, -18246, -15960, -12598, -14486, -28329, -40490, -31319, -7952, 657, -15831, -35487, -36772, -24243, -12673, -5511, -2311, -9437, -25482, -30192, -9126, 19530, 24844, 5447, -9852, -2557, 16510, 30895, 38336, 39908, 31520, 18804, 21432, 45866, 68469, 64470, 42914, 32951, 43357, 57234, 62299, 62881, 61428, 52203, 39608, 40547, 57687, 69331, 59531, 42018, 38357, 46595, 50475, 48395, 50949, 56230, 51666, 39761, 38568, 52410, 63591, 60569, 54303, 56340, 59885, 56962, 57159};
// always_comb correct_outputs = '{-680344, -1249027, -729189, 1604747, 5510102, 9517597, 11225695, 8257649, -193474, -12036352, -22348746, -25225238, -16561402, 3491148, 29339678, 50756621, 56169119, 37863337, -3036453, -54530355, -96273242, -106458679, -71194131, 6905391, 105038314, 184675544, 204221742, 136129330, -17532302, -217019524, -388544939, -440467321, -288384022, 118584483, 779191628, 1635563348, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2119050508, 1961578198, 1825613808, 1711726412, 1618520094, 1543913620, 1486144420, 1443869537, 1415644487, 1399583439, 1393463392, 1395334482, 1401729440, 1409349257, 1415045527, 1415850343, 1408712506, 1390536666, 1358577801, 1310619698, 1244769489, 1159378250, 1053322259, 926173231, 777959263, 608969735, 420003136, 212650657, -10913061, -248349975, -497174709, -754468102, -1016886292, -1281003119, -1543457205, -1800804872, -2049565754, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116424109, -1966200130, -1833456980, -1719204103, -1623656724, -1546414429, -1486748438, -1443526511, -1415026426, -1399085387, -1393370079, -1395295928, -1401790068, -1409464270, -1415100177, -1415786123, -1408603216, -1390497512, -1358629108, -1310688480, -1244798133, -1159370150, -1053293395, -926128433, -777925344, -608988455, -420066199, -212691504, 10934638, 248397668, 497197646, 754467482, 1016883018, 1280984437, 1543410748, 1800774184, 2049604907, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2116432099, 1966254228, 1833495929, 1719199916, 1623634864, 1546392840, 1486718012, 1443502820, 1415054996, 1399162709, 1393414651, 1395245950, 1401693470, 1409422554, 1415147310, 1415868176, 1408654856, 1390489290, 1358560455, 1310596159, 1244764317, 1159451978, 1053428891, 926175129, 777824466, 608843488, 420023277, 212780111, -10808148, -248337736, -497242634, -754585812, -1016987672, -1280976052, -1543274751, -1800632613, -2049607436, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116288505, -1966208814, -1833573049, -1719323701, -1623710967, -1546362187, -1486591395, -1443380596, -1415061729, -1399309517, -1393558099, -1395236836, -1401547290, -1409293513, -1415149926, -1415976828, -1408766703, -1390523934, -1358496187, -1310475479, -1244686307, -1159499955, -1053567883, -926264615, -777772732, -608714815, -419953035, -212818149, 10723054, 248279976, 497238088, 754630761, 1017059437, 1281019096, 1543239093, 1800546637, 2049562238};

// module fir #(clk, rst, ena, sample, out);
fir UUT(.clk(clk), .rst(rst), .ena(shift_ena), .sample(next_sample), .out(out));

// Some behavioural comb. logic that computes correct values.

// toggle every two clock cycles
logic toggle;
always_ff @(posedge clk) begin
    toggle <= ~toggle;
    if (toggle) begin
        counter <= counter + 1;
        #1 print_io();
        assert(out === correct_out) else begin
        // $display("  ERROR: mux out should be %b, is %b", out, correct_out);
        errors = errors + 1;
  end
    end else begin
        counter <= counter;
    end
end

always_comb begin : simulated_output
  next_sample <= samples[counter];
  correct_out = correct_outputs[counter];
end

task print_io;
  $display("%b | %b (%b)", counter, next_sample, correct_out);
endtask

initial begin
  # 1;
  if (errors !== 0) begin
    $display("---------------------------------------------------------------");
    $display("-- FAILURE                                                   --");
    $display("---------------------------------------------------------------");
    $display(" %d failures found, try again!", errors);
  end else begin
    $display("---------------------------------------------------------------");
    $display("-- SUCCESS                                                   --");
    $display("---------------------------------------------------------------");
  end
  $finish;
end

always #(10) clk = ~clk;

endmodule
