`timescale 1ns/1ps
`default_nettype none

module test_fir;
int errors = 0;

// PASTE COPIED CODE BELOW

logic rst;
logic clk;
logic shift_ena;
logic [15:0] next_sample;
logic [38:0] out;
logic signed [39:0] diff;

integer counter;
logic [38:0] correct_out;

logic [6399:0] packed_samples;
always_comb packed_samples = {16'sd3572, 16'sd3560, 16'sd3742, 16'sd3521, 16'sd3393, 16'sd3785, 16'sd3974, 16'sd3275, 16'sd2410, 16'sd2485, 16'sd3229, 16'sd3514, 16'sd3184, 16'sd3024, 16'sd3154, 16'sd2912, 16'sd2397, 16'sd2626, 16'sd3720, 16'sd4333, 16'sd3605, 16'sd2534, 16'sd2475, 16'sd3262, 16'sd3839, 16'sd3930, 16'sd3893, 16'sd3577, 16'sd2709, 16'sd2059, 16'sd2682, 16'sd4029, 16'sd4279, 16'sd2866, 16'sd1339, 16'sd1175, 16'sd1970, 16'sd2494, 16'sd2396, 16'sd1930, 16'sd1031, -16'sd159, -16'sd615, 16'sd340, 16'sd1552, 16'sd1220, -16'sd570, -16'sd1887, -16'sd1592, -16'sd589, -16'sd144, -16'sd344, -16'sd792, -16'sd1515, -16'sd2298, -16'sd2217, -16'sd989, 16'sd41, -16'sd497, -16'sd1957, -16'sd2530, -16'sd1770, -16'sd905, -16'sd787, -16'sd997, -16'sd1140, -16'sd1546, -16'sd2175, -16'sd2165, -16'sd1281, -16'sd693, -16'sd1345, -16'sd2458, -16'sd2741, -16'sd2329, -16'sd2259, -16'sd2637, -16'sd2717, -16'sd2543, -16'sd2968, -16'sd3972, -16'sd4411, -16'sd3850, -16'sd3325, -16'sd3692, -16'sd4395, -16'sd4641, -16'sd4698, -16'sd5030, -16'sd5129, -16'sd4436, -16'sd3744, -16'sd4231, -16'sd5472, -16'sd5840, -16'sd4863, -16'sd3789, -16'sd3638, -16'sd4031, -16'sd4328, -16'sd4586, -16'sd4749, -16'sd4159, -16'sd2823, -16'sd2125, -16'sd3060, -16'sd4514, -16'sd4595, -16'sd3221, -16'sd2044, -16'sd2076, -16'sd2772, -16'sd3392, -16'sd3835, -16'sd3882, -16'sd3064, -16'sd1874, -16'sd1808, -16'sd3303, -16'sd4726, -16'sd4431, -16'sd2985, -16'sd2202, -16'sd2662, -16'sd3462, -16'sd3926, -16'sd4141, -16'sd3972, -16'sd3075, -16'sd2062, -16'sd2194, -16'sd3448, -16'sd4167, -16'sd3312, -16'sd1909, -16'sd1436, -16'sd1799, -16'sd1988, -16'sd1820, -16'sd1756, -16'sd1586, -16'sd762, 16'sd233, 16'sd296, -16'sd474, -16'sd742, 16'sd31, 16'sd853, 16'sd931, 16'sd817, 16'sd1131, 16'sd1345, 16'sd888, 16'sd456, 16'sd982, 16'sd1955, 16'sd2103, 16'sd1368, 16'sd854, 16'sd1000, 16'sd1191, 16'sd1191, 16'sd1524, 16'sd2102, 16'sd1928, 16'sd814, 16'sd147, 16'sd976, 16'sd2359, 16'sd2694, 16'sd1928, 16'sd1261, 16'sd1263, 16'sd1590, 16'sd2151, 16'sd3101, 16'sd3791, 16'sd3249, 16'sd1959, 16'sd1729, 16'sd3225, 16'sd4885, 16'sd5048, 16'sd4057, 16'sd3356, 16'sd3470, 16'sd3988, 16'sd4732, 16'sd5602, 16'sd5812, 16'sd4745, 16'sd3392, 16'sd3474, 16'sd5004, 16'sd6093, 16'sd5522, 16'sd4206, 16'sd3561, 16'sd3687, 16'sd3972, 16'sd4329, 16'sd4756, 16'sd4572, 16'sd3397, 16'sd2298, 16'sd2596, 16'sd3838, 16'sd4323, 16'sd3530, 16'sd2646, 16'sd2564, 16'sd2805, 16'sd2824, 16'sd2995, 16'sd3543, 16'sd3707, 16'sd2991, 16'sd2289, 16'sd2642, 16'sd3565, 16'sd3841, 16'sd3434, 16'sd3277, 16'sd3506, 16'sd3366, 16'sd2856, 16'sd2944, 16'sd3800, 16'sd4226, 16'sd3482, 16'sd2478, 16'sd2329, 16'sd2757, 16'sd2899, 16'sd2765, 16'sd2760, 16'sd2501, 16'sd1486, 16'sd476, 16'sd714, 16'sd1862, 16'sd2177, 16'sd970, -16'sd476, -16'sd851, -16'sd407, -16'sd12, 16'sd160, 16'sd143, -16'sd515, -16'sd1803, -16'sd2463, -16'sd1503, 16'sd29, 16'sd181, -16'sd1239, -16'sd2495, -16'sd2381, -16'sd1488, -16'sd812, -16'sd523, -16'sd610, -16'sd1370, -16'sd2452, -16'sd2571, -16'sd1246, 16'sd50, -16'sd321, -16'sd1882, -16'sd2785, -16'sd2372, -16'sd1644, -16'sd1418, -16'sd1508, -16'sd1790, -16'sd2594, -16'sd3590, -16'sd3680, -16'sd2696, -16'sd2052, -16'sd2824, -16'sd4153, -16'sd4598, -16'sd4196, -16'sd3995, -16'sd4204, -16'sd4211, -16'sd4084, -16'sd4525, -16'sd5351, -16'sd5462, -16'sd4641, -16'sd4036, -16'sd4369, -16'sd4892, -16'sd4805, -16'sd4535, -16'sd4679, -16'sd4717, -16'sd3990, -16'sd3175, -16'sd3410, -16'sd4361, -16'sd4601, -16'sd3753, -16'sd2898, -16'sd2775, -16'sd2950, -16'sd3038, -16'sd3369, -16'sd3873, -16'sd3630, -16'sd2423, -16'sd1634, -16'sd2441, -16'sd3953, -16'sd4367, -16'sd3437, -16'sd2494, -16'sd2392, -16'sd2796, -16'sd3352, -16'sd4088, -16'sd4512, -16'sd3790, -16'sd2336, -16'sd1878, -16'sd3147, -16'sd4621, -16'sd4517, -16'sd3123, -16'sd2053, -16'sd1983, -16'sd2360, -16'sd2769, -16'sd3164, -16'sd3030, -16'sd1821, -16'sd323, -16'sd127, -16'sd1353, -16'sd2224, -16'sd1475, 16'sd17, 16'sd748, 16'sd604, 16'sd377, 16'sd248, 16'sd17, 16'sd130, 16'sd1074, 16'sd2093, 16'sd1934, 16'sd816, 16'sd283, 16'sd945, 16'sd1730, 16'sd1731, 16'sd1441, 16'sd1503, 16'sd1503, 16'sd989, 16'sd634, 16'sd1188, 16'sd2026, 16'sd2001, 16'sd1269, 16'sd961, 16'sd1322, 16'sd1568, 16'sd1511, 16'sd1844, 16'sd2586, 16'sd2706, 16'sd1887, 16'sd1369, 16'sd2157, 16'sd3455, 16'sd3897, 16'sd3482, 16'sd3158, 16'sd3203, 16'sd3281, 16'sd3604, 16'sd4577, 16'sd5499, 16'sd5135, 16'sd3759, 16'sd3176, 16'sd4251, 16'sd5683, 16'sd5913, 16'sd5083, 16'sd4285, 16'sd3923, 16'sd3867, 16'sd4328, 16'sd5285, 16'sd5660, 16'sd4512};
logic [15:0] samples[0:399];
always_comb begin 
samples[0] = packed_samples[15:0]; samples[1] = packed_samples[31:16]; samples[2] = packed_samples[47:32]; samples[3] = packed_samples[63:48]; samples[4] = packed_samples[79:64]; samples[5] = packed_samples[95:80]; samples[6] = packed_samples[111:96]; samples[7] = packed_samples[127:112]; samples[8] = packed_samples[143:128]; samples[9] = packed_samples[159:144]; samples[10] = packed_samples[175:160]; samples[11] = packed_samples[191:176]; samples[12] = packed_samples[207:192]; samples[13] = packed_samples[223:208]; samples[14] = packed_samples[239:224]; samples[15] = packed_samples[255:240]; samples[16] = packed_samples[271:256]; samples[17] = packed_samples[287:272]; samples[18] = packed_samples[303:288]; samples[19] = packed_samples[319:304]; samples[20] = packed_samples[335:320]; samples[21] = packed_samples[351:336]; samples[22] = packed_samples[367:352]; samples[23] = packed_samples[383:368]; samples[24] = packed_samples[399:384]; samples[25] = packed_samples[415:400]; samples[26] = packed_samples[431:416]; samples[27] = packed_samples[447:432]; samples[28] = packed_samples[463:448]; samples[29] = packed_samples[479:464]; samples[30] = packed_samples[495:480]; samples[31] = packed_samples[511:496]; samples[32] = packed_samples[527:512]; samples[33] = packed_samples[543:528]; samples[34] = packed_samples[559:544]; samples[35] = packed_samples[575:560]; samples[36] = packed_samples[591:576]; samples[37] = packed_samples[607:592]; samples[38] = packed_samples[623:608]; samples[39] = packed_samples[639:624]; samples[40] = packed_samples[655:640]; samples[41] = packed_samples[671:656]; samples[42] = packed_samples[687:672]; samples[43] = packed_samples[703:688]; samples[44] = packed_samples[719:704]; samples[45] = packed_samples[735:720]; samples[46] = packed_samples[751:736]; samples[47] = packed_samples[767:752]; samples[48] = packed_samples[783:768]; samples[49] = packed_samples[799:784]; samples[50] = packed_samples[815:800]; samples[51] = packed_samples[831:816]; samples[52] = packed_samples[847:832]; samples[53] = packed_samples[863:848]; samples[54] = packed_samples[879:864]; samples[55] = packed_samples[895:880]; samples[56] = packed_samples[911:896]; samples[57] = packed_samples[927:912]; samples[58] = packed_samples[943:928]; samples[59] = packed_samples[959:944]; samples[60] = packed_samples[975:960]; samples[61] = packed_samples[991:976]; samples[62] = packed_samples[1007:992]; samples[63] = packed_samples[1023:1008]; samples[64] = packed_samples[1039:1024]; samples[65] = packed_samples[1055:1040]; samples[66] = packed_samples[1071:1056]; samples[67] = packed_samples[1087:1072]; samples[68] = packed_samples[1103:1088]; samples[69] = packed_samples[1119:1104]; samples[70] = packed_samples[1135:1120]; samples[71] = packed_samples[1151:1136]; samples[72] = packed_samples[1167:1152]; samples[73] = packed_samples[1183:1168]; samples[74] = packed_samples[1199:1184]; samples[75] = packed_samples[1215:1200]; samples[76] = packed_samples[1231:1216]; samples[77] = packed_samples[1247:1232]; samples[78] = packed_samples[1263:1248]; samples[79] = packed_samples[1279:1264]; samples[80] = packed_samples[1295:1280]; samples[81] = packed_samples[1311:1296]; samples[82] = packed_samples[1327:1312]; samples[83] = packed_samples[1343:1328]; samples[84] = packed_samples[1359:1344]; samples[85] = packed_samples[1375:1360]; samples[86] = packed_samples[1391:1376]; samples[87] = packed_samples[1407:1392]; samples[88] = packed_samples[1423:1408]; samples[89] = packed_samples[1439:1424]; samples[90] = packed_samples[1455:1440]; samples[91] = packed_samples[1471:1456]; samples[92] = packed_samples[1487:1472]; samples[93] = packed_samples[1503:1488]; samples[94] = packed_samples[1519:1504]; samples[95] = packed_samples[1535:1520]; samples[96] = packed_samples[1551:1536]; samples[97] = packed_samples[1567:1552]; samples[98] = packed_samples[1583:1568]; samples[99] = packed_samples[1599:1584]; samples[100] = packed_samples[1615:1600]; samples[101] = packed_samples[1631:1616]; samples[102] = packed_samples[1647:1632]; samples[103] = packed_samples[1663:1648]; samples[104] = packed_samples[1679:1664]; samples[105] = packed_samples[1695:1680]; samples[106] = packed_samples[1711:1696]; samples[107] = packed_samples[1727:1712]; samples[108] = packed_samples[1743:1728]; samples[109] = packed_samples[1759:1744]; samples[110] = packed_samples[1775:1760]; samples[111] = packed_samples[1791:1776]; samples[112] = packed_samples[1807:1792]; samples[113] = packed_samples[1823:1808]; samples[114] = packed_samples[1839:1824]; samples[115] = packed_samples[1855:1840]; samples[116] = packed_samples[1871:1856]; samples[117] = packed_samples[1887:1872]; samples[118] = packed_samples[1903:1888]; samples[119] = packed_samples[1919:1904]; samples[120] = packed_samples[1935:1920]; samples[121] = packed_samples[1951:1936]; samples[122] = packed_samples[1967:1952]; samples[123] = packed_samples[1983:1968]; samples[124] = packed_samples[1999:1984]; samples[125] = packed_samples[2015:2000]; samples[126] = packed_samples[2031:2016]; samples[127] = packed_samples[2047:2032]; samples[128] = packed_samples[2063:2048]; samples[129] = packed_samples[2079:2064]; samples[130] = packed_samples[2095:2080]; samples[131] = packed_samples[2111:2096]; samples[132] = packed_samples[2127:2112]; samples[133] = packed_samples[2143:2128]; samples[134] = packed_samples[2159:2144]; samples[135] = packed_samples[2175:2160]; samples[136] = packed_samples[2191:2176]; samples[137] = packed_samples[2207:2192]; samples[138] = packed_samples[2223:2208]; samples[139] = packed_samples[2239:2224]; samples[140] = packed_samples[2255:2240]; samples[141] = packed_samples[2271:2256]; samples[142] = packed_samples[2287:2272]; samples[143] = packed_samples[2303:2288]; samples[144] = packed_samples[2319:2304]; samples[145] = packed_samples[2335:2320]; samples[146] = packed_samples[2351:2336]; samples[147] = packed_samples[2367:2352]; samples[148] = packed_samples[2383:2368]; samples[149] = packed_samples[2399:2384]; samples[150] = packed_samples[2415:2400]; samples[151] = packed_samples[2431:2416]; samples[152] = packed_samples[2447:2432]; samples[153] = packed_samples[2463:2448]; samples[154] = packed_samples[2479:2464]; samples[155] = packed_samples[2495:2480]; samples[156] = packed_samples[2511:2496]; samples[157] = packed_samples[2527:2512]; samples[158] = packed_samples[2543:2528]; samples[159] = packed_samples[2559:2544]; samples[160] = packed_samples[2575:2560]; samples[161] = packed_samples[2591:2576]; samples[162] = packed_samples[2607:2592]; samples[163] = packed_samples[2623:2608]; samples[164] = packed_samples[2639:2624]; samples[165] = packed_samples[2655:2640]; samples[166] = packed_samples[2671:2656]; samples[167] = packed_samples[2687:2672]; samples[168] = packed_samples[2703:2688]; samples[169] = packed_samples[2719:2704]; samples[170] = packed_samples[2735:2720]; samples[171] = packed_samples[2751:2736]; samples[172] = packed_samples[2767:2752]; samples[173] = packed_samples[2783:2768]; samples[174] = packed_samples[2799:2784]; samples[175] = packed_samples[2815:2800]; samples[176] = packed_samples[2831:2816]; samples[177] = packed_samples[2847:2832]; samples[178] = packed_samples[2863:2848]; samples[179] = packed_samples[2879:2864]; samples[180] = packed_samples[2895:2880]; samples[181] = packed_samples[2911:2896]; samples[182] = packed_samples[2927:2912]; samples[183] = packed_samples[2943:2928]; samples[184] = packed_samples[2959:2944]; samples[185] = packed_samples[2975:2960]; samples[186] = packed_samples[2991:2976]; samples[187] = packed_samples[3007:2992]; samples[188] = packed_samples[3023:3008]; samples[189] = packed_samples[3039:3024]; samples[190] = packed_samples[3055:3040]; samples[191] = packed_samples[3071:3056]; samples[192] = packed_samples[3087:3072]; samples[193] = packed_samples[3103:3088]; samples[194] = packed_samples[3119:3104]; samples[195] = packed_samples[3135:3120]; samples[196] = packed_samples[3151:3136]; samples[197] = packed_samples[3167:3152]; samples[198] = packed_samples[3183:3168]; samples[199] = packed_samples[3199:3184]; samples[200] = packed_samples[3215:3200]; samples[201] = packed_samples[3231:3216]; samples[202] = packed_samples[3247:3232]; samples[203] = packed_samples[3263:3248]; samples[204] = packed_samples[3279:3264]; samples[205] = packed_samples[3295:3280]; samples[206] = packed_samples[3311:3296]; samples[207] = packed_samples[3327:3312]; samples[208] = packed_samples[3343:3328]; samples[209] = packed_samples[3359:3344]; samples[210] = packed_samples[3375:3360]; samples[211] = packed_samples[3391:3376]; samples[212] = packed_samples[3407:3392]; samples[213] = packed_samples[3423:3408]; samples[214] = packed_samples[3439:3424]; samples[215] = packed_samples[3455:3440]; samples[216] = packed_samples[3471:3456]; samples[217] = packed_samples[3487:3472]; samples[218] = packed_samples[3503:3488]; samples[219] = packed_samples[3519:3504]; samples[220] = packed_samples[3535:3520]; samples[221] = packed_samples[3551:3536]; samples[222] = packed_samples[3567:3552]; samples[223] = packed_samples[3583:3568]; samples[224] = packed_samples[3599:3584]; samples[225] = packed_samples[3615:3600]; samples[226] = packed_samples[3631:3616]; samples[227] = packed_samples[3647:3632]; samples[228] = packed_samples[3663:3648]; samples[229] = packed_samples[3679:3664]; samples[230] = packed_samples[3695:3680]; samples[231] = packed_samples[3711:3696]; samples[232] = packed_samples[3727:3712]; samples[233] = packed_samples[3743:3728]; samples[234] = packed_samples[3759:3744]; samples[235] = packed_samples[3775:3760]; samples[236] = packed_samples[3791:3776]; samples[237] = packed_samples[3807:3792]; samples[238] = packed_samples[3823:3808]; samples[239] = packed_samples[3839:3824]; samples[240] = packed_samples[3855:3840]; samples[241] = packed_samples[3871:3856]; samples[242] = packed_samples[3887:3872]; samples[243] = packed_samples[3903:3888]; samples[244] = packed_samples[3919:3904]; samples[245] = packed_samples[3935:3920]; samples[246] = packed_samples[3951:3936]; samples[247] = packed_samples[3967:3952]; samples[248] = packed_samples[3983:3968]; samples[249] = packed_samples[3999:3984]; samples[250] = packed_samples[4015:4000]; samples[251] = packed_samples[4031:4016]; samples[252] = packed_samples[4047:4032]; samples[253] = packed_samples[4063:4048]; samples[254] = packed_samples[4079:4064]; samples[255] = packed_samples[4095:4080]; samples[256] = packed_samples[4111:4096]; samples[257] = packed_samples[4127:4112]; samples[258] = packed_samples[4143:4128]; samples[259] = packed_samples[4159:4144]; samples[260] = packed_samples[4175:4160]; samples[261] = packed_samples[4191:4176]; samples[262] = packed_samples[4207:4192]; samples[263] = packed_samples[4223:4208]; samples[264] = packed_samples[4239:4224]; samples[265] = packed_samples[4255:4240]; samples[266] = packed_samples[4271:4256]; samples[267] = packed_samples[4287:4272]; samples[268] = packed_samples[4303:4288]; samples[269] = packed_samples[4319:4304]; samples[270] = packed_samples[4335:4320]; samples[271] = packed_samples[4351:4336]; samples[272] = packed_samples[4367:4352]; samples[273] = packed_samples[4383:4368]; samples[274] = packed_samples[4399:4384]; samples[275] = packed_samples[4415:4400]; samples[276] = packed_samples[4431:4416]; samples[277] = packed_samples[4447:4432]; samples[278] = packed_samples[4463:4448]; samples[279] = packed_samples[4479:4464]; samples[280] = packed_samples[4495:4480]; samples[281] = packed_samples[4511:4496]; samples[282] = packed_samples[4527:4512]; samples[283] = packed_samples[4543:4528]; samples[284] = packed_samples[4559:4544]; samples[285] = packed_samples[4575:4560]; samples[286] = packed_samples[4591:4576]; samples[287] = packed_samples[4607:4592]; samples[288] = packed_samples[4623:4608]; samples[289] = packed_samples[4639:4624]; samples[290] = packed_samples[4655:4640]; samples[291] = packed_samples[4671:4656]; samples[292] = packed_samples[4687:4672]; samples[293] = packed_samples[4703:4688]; samples[294] = packed_samples[4719:4704]; samples[295] = packed_samples[4735:4720]; samples[296] = packed_samples[4751:4736]; samples[297] = packed_samples[4767:4752]; samples[298] = packed_samples[4783:4768]; samples[299] = packed_samples[4799:4784]; samples[300] = packed_samples[4815:4800]; samples[301] = packed_samples[4831:4816]; samples[302] = packed_samples[4847:4832]; samples[303] = packed_samples[4863:4848]; samples[304] = packed_samples[4879:4864]; samples[305] = packed_samples[4895:4880]; samples[306] = packed_samples[4911:4896]; samples[307] = packed_samples[4927:4912]; samples[308] = packed_samples[4943:4928]; samples[309] = packed_samples[4959:4944]; samples[310] = packed_samples[4975:4960]; samples[311] = packed_samples[4991:4976]; samples[312] = packed_samples[5007:4992]; samples[313] = packed_samples[5023:5008]; samples[314] = packed_samples[5039:5024]; samples[315] = packed_samples[5055:5040]; samples[316] = packed_samples[5071:5056]; samples[317] = packed_samples[5087:5072]; samples[318] = packed_samples[5103:5088]; samples[319] = packed_samples[5119:5104]; samples[320] = packed_samples[5135:5120]; samples[321] = packed_samples[5151:5136]; samples[322] = packed_samples[5167:5152]; samples[323] = packed_samples[5183:5168]; samples[324] = packed_samples[5199:5184]; samples[325] = packed_samples[5215:5200]; samples[326] = packed_samples[5231:5216]; samples[327] = packed_samples[5247:5232]; samples[328] = packed_samples[5263:5248]; samples[329] = packed_samples[5279:5264]; samples[330] = packed_samples[5295:5280]; samples[331] = packed_samples[5311:5296]; samples[332] = packed_samples[5327:5312]; samples[333] = packed_samples[5343:5328]; samples[334] = packed_samples[5359:5344]; samples[335] = packed_samples[5375:5360]; samples[336] = packed_samples[5391:5376]; samples[337] = packed_samples[5407:5392]; samples[338] = packed_samples[5423:5408]; samples[339] = packed_samples[5439:5424]; samples[340] = packed_samples[5455:5440]; samples[341] = packed_samples[5471:5456]; samples[342] = packed_samples[5487:5472]; samples[343] = packed_samples[5503:5488]; samples[344] = packed_samples[5519:5504]; samples[345] = packed_samples[5535:5520]; samples[346] = packed_samples[5551:5536]; samples[347] = packed_samples[5567:5552]; samples[348] = packed_samples[5583:5568]; samples[349] = packed_samples[5599:5584]; samples[350] = packed_samples[5615:5600]; samples[351] = packed_samples[5631:5616]; samples[352] = packed_samples[5647:5632]; samples[353] = packed_samples[5663:5648]; samples[354] = packed_samples[5679:5664]; samples[355] = packed_samples[5695:5680]; samples[356] = packed_samples[5711:5696]; samples[357] = packed_samples[5727:5712]; samples[358] = packed_samples[5743:5728]; samples[359] = packed_samples[5759:5744]; samples[360] = packed_samples[5775:5760]; samples[361] = packed_samples[5791:5776]; samples[362] = packed_samples[5807:5792]; samples[363] = packed_samples[5823:5808]; samples[364] = packed_samples[5839:5824]; samples[365] = packed_samples[5855:5840]; samples[366] = packed_samples[5871:5856]; samples[367] = packed_samples[5887:5872]; samples[368] = packed_samples[5903:5888]; samples[369] = packed_samples[5919:5904]; samples[370] = packed_samples[5935:5920]; samples[371] = packed_samples[5951:5936]; samples[372] = packed_samples[5967:5952]; samples[373] = packed_samples[5983:5968]; samples[374] = packed_samples[5999:5984]; samples[375] = packed_samples[6015:6000]; samples[376] = packed_samples[6031:6016]; samples[377] = packed_samples[6047:6032]; samples[378] = packed_samples[6063:6048]; samples[379] = packed_samples[6079:6064]; samples[380] = packed_samples[6095:6080]; samples[381] = packed_samples[6111:6096]; samples[382] = packed_samples[6127:6112]; samples[383] = packed_samples[6143:6128]; samples[384] = packed_samples[6159:6144]; samples[385] = packed_samples[6175:6160]; samples[386] = packed_samples[6191:6176]; samples[387] = packed_samples[6207:6192]; samples[388] = packed_samples[6223:6208]; samples[389] = packed_samples[6239:6224]; samples[390] = packed_samples[6255:6240]; samples[391] = packed_samples[6271:6256]; samples[392] = packed_samples[6287:6272]; samples[393] = packed_samples[6303:6288]; samples[394] = packed_samples[6319:6304]; samples[395] = packed_samples[6335:6320]; samples[396] = packed_samples[6351:6336]; samples[397] = packed_samples[6367:6352]; samples[398] = packed_samples[6383:6368]; samples[399] = packed_samples[6399:6384]; 
end

logic [15599:0] packed_outputs;
always_comb packed_outputs = {39'sd128097639, 39'sd112534164, 39'sd96452443, 39'sd80063693, 39'sd63566214, 39'sd47164422, 39'sd31077380, 39'sd15517498, 39'sd670190, -39'sd13301134, -39'sd26247064, -39'sd38044675, -39'sd48610795, -39'sd57891538, -39'sd65847992, -39'sd72468747, -39'sd77792894, -39'sd81904717, -39'sd84906011, -39'sd86907745, -39'sd88047918, -39'sd88498551, -39'sd88446870, -39'sd88080844, -39'sd87596705, -39'sd87202302, -39'sd87097381, -39'sd87456844, -39'sd88441358, -39'sd90211287, -39'sd92911962, -39'sd96647636, -39'sd101481935, -39'sd107457731, -39'sd114598315, -39'sd122888050, -39'sd132268031, -39'sd142654464, -39'sd153946632, -39'sd166011953, -39'sd178679716, -39'sd191761676, -39'sd205070277, -39'sd218409732, -39'sd231564136, -39'sd244312183, -39'sd256450188, -39'sd267790415, -39'sd278146699, -39'sd287342694, -39'sd295236989, -39'sd301727435, -39'sd306732167, -39'sd310184618, -39'sd312053745, -39'sd312355741, -39'sd311139318, -39'sd308472914, -39'sd304454994, -39'sd299222963, -39'sd292936946, -39'sd285761315, -39'sd277873180, -39'sd269478628, -39'sd260800464, -39'sd252048280, -39'sd243411515, -39'sd235076754, -39'sd227231297, -39'sd220042816, -39'sd213646959, -39'sd208156616, -39'sd203665113, -39'sd200228892, -39'sd197858268, -39'sd196535557, -39'sd196231351, -39'sd196889839, -39'sd198406883, -39'sd200638808, -39'sd203430041, -39'sd206619771, -39'sd210027639, -39'sd213453300, -39'sd216695211, -39'sd219558124, -39'sd221842718, -39'sd223348224, -39'sd223897496, -39'sd223350418, -39'sd221587006, -39'sd218492702, -39'sd213975319, -39'sd207989423, -39'sd200532358, -39'sd191624804, -39'sd181311170, -39'sd169674630, -39'sd156834213, -39'sd142925901, -39'sd128100464, -39'sd112539538, -39'sd96454671, -39'sd80061003, -39'sd63561729, -39'sd47161613, -39'sd31077664, -39'sd15521108, -39'sd675509, 39'sd13298756, 39'sd26251454, 39'sd38052718, 39'sd48614029, 39'sd57885945, 39'sd65839305, 39'sd72465748, 39'sd77797769, 39'sd81912259, 39'sd84910028, 39'sd86905580, 39'sd88040928, 39'sd88491761, 39'sd88446706, 39'sd88088909, 39'sd87605841, 39'sd87202871, 39'sd87088415, 39'sd87447669, 39'sd88440937, 39'sd90218926, 39'sd92919875, 39'sd96649552, 39'sd101477179, 39'sd107449994, 39'sd114593495, 39'sd122890889, 39'sd132277006, 39'sd142661137, 39'sd153943860, 39'sd166002527, 39'sd178673537, 39'sd191764347, 39'sd205077796, 39'sd218414693, 39'sd231563444, 39'sd244307570, 39'sd256444999, 39'sd267788211, 39'sd278149849, 39'sd287349151, 39'sd295240492, 39'sd301724147, 39'sd306725803, 39'sd310182015, 39'sd312056549, 39'sd312359715, 39'sd311140910, 39'sd308472523, 39'sd304453781, 39'sd299220742, 39'sd292934597, 39'sd285761539, 39'sd277876564, 39'sd269481695, 39'sd260800032, 39'sd252045568, 39'sd243409606, 39'sd235076244, 39'sd227231284, 39'sd220044049, 39'sd213650203, 39'sd208159084, 39'sd203662908, 39'sd200223227, 39'sd197855271, 39'sd196538682, 39'sd196237155, 39'sd196892688, 39'sd198405011, 39'sd200634277, 39'sd203425776, 39'sd206618747, 39'sd210031893, 39'sd213460461, 39'sd216698264, 39'sd219552675, 39'sd221833605, 39'sd223345036, 39'sd223903475, 39'sd223359123, 39'sd221590236, 39'sd218488532, 39'sd213967869, 39'sd207984319, 39'sd200533614, 39'sd191632385, 39'sd181319162, 39'sd169674919, 39'sd156825375, 39'sd142916531, 39'sd128100306, 39'sd112548386, 39'sd96463171, 39'sd80061527, 39'sd63555188, 39'sd47154217, 39'sd31074852, 39'sd15524854, 39'sd683414, -39'sd13293219, -39'sd26254137, -39'sd38061778, -39'sd48620334, -39'sd57883027, -39'sd65830837, -39'sd72460634, -39'sd77799883, -39'sd81918030, -39'sd84914319, -39'sd86906094, -39'sd88037701, -39'sd88486632, -39'sd88443761, -39'sd88091516, -39'sd87611879, -39'sd87205995, -39'sd87085629, -39'sd87442836, -39'sd88439151, -39'sd90220406, -39'sd92921777, -39'sd96650901, -39'sd101478545, -39'sd107450256, -39'sd114591061, -39'sd122887508, -39'sd132276506, -39'sd142664116, -39'sd153946888, -39'sd166003041, -39'sd178672327, -39'sd191762638, -39'sd205075487, -39'sd218412924, -39'sd231565155, -39'sd244312779, -39'sd256448454, -39'sd267785290, -39'sd278143154, -39'sd287345754, -39'sd295243489, -39'sd301730036, -39'sd306729512, -39'sd310181269, -39'sd312051824, -39'sd312353787, -39'sd311138802, -39'sd308477668, -39'sd304462477, -39'sd299224019, -39'sd292928282, -39'sd285751967, -39'sd277873515, -39'sd269487528, -39'sd260808448, -39'sd252049317, -39'sd243406407, -39'sd235068734, -39'sd227224990, -39'sd220044654, -39'sd213658473, -39'sd208167845, -39'sd203662985, -39'sd200214003, -39'sd197846262, -39'sd196538839, -39'sd196245284, -39'sd196900328, -39'sd198406014, -39'sd200629046, -39'sd203418701, -39'sd206614984, -39'sd210034891, -39'sd213468534, -39'sd216704066, -39'sd219549960, -39'sd221824950, -39'sd223339560, -39'sd223906260, -39'sd223366079, -39'sd221594301, -39'sd218487402, -39'sd213963922, -39'sd207980417, -39'sd200531898, -39'sd191634533, -39'sd181324185, -39'sd169678164, -39'sd156823220, -39'sd142911400, -39'sd128097859, -39'sd112550304, -39'sd96466075, -39'sd80062694, -39'sd63555393, -39'sd47154256, -39'sd31073419, -39'sd15521873, -39'sd682066, 39'sd13290666, 39'sd26250196, 39'sd38060608, 39'sd48622453, 39'sd57885826, 39'sd65832641, 39'sd72461140, 39'sd77798093, 39'sd81913731, 39'sd84911112, 39'sd86908541, 39'sd88044531, 39'sd88490646, 39'sd88440345, 39'sd88084328, 39'sd87608090, 39'sd87208405, 39'sd87091462, 39'sd87473964, 39'sd88477780, 39'sd90241846, 39'sd92884026, 39'sd96494601, 39'sd101157505, 39'sd106982900, 39'sd114100863, 39'sd122598637, 39'sd132440656, 39'sd143422031, 39'sd155180921, 39'sd167280139, 39'sd179354210, 39'sd191269907, 39'sd203200364, 39'sd215538792, 39'sd228671271, 39'sd242702472, 39'sd257240305, 39'sd271334444, 39'sd283648215, 39'sd292875810, 39'sd298283909, 39'sd300146685, 39'sd299848987, 39'sd299543926, 39'sd301400966, 39'sd306638457, 39'sd314678486, 39'sd322806906, 39'sd326581852, 39'sd320952131, 39'sd301774473, 39'sd267267712, 39'sd218927163, 39'sd161541829, 39'sd102222709, 39'sd48699476, 39'sd7411530, -39'sd18024001, -39'sd27529207, -39'sd24284058, -39'sd13563720, -39'sd1095768, 39'sd8508083, 39'sd12763858, 39'sd11542221, 39'sd6564894, 39'sd431586, -39'sd4449633, -39'sd6653667, -39'sd6017077, -39'sd3408147, -39'sd189778, 39'sd2366458, 39'sd3510569, 39'sd3172288, 39'sd1833729, 39'sd218196, -39'sd1035087, -39'sd1576577, -39'sd1396796, -39'sd752272, -39'sd12092, 39'sd516103, 39'sd701605, 39'sd594849, 39'sd344381, 39'sd100296, -39'sd45574, -39'sd78064, -39'sd42521};
logic [38:0] correct_outputs[0:399];
always_comb begin
correct_outputs[0] = packed_outputs[38:0]; correct_outputs[1] = packed_outputs[77:39]; correct_outputs[2] = packed_outputs[116:78]; correct_outputs[3] = packed_outputs[155:117]; correct_outputs[4] = packed_outputs[194:156]; correct_outputs[5] = packed_outputs[233:195]; correct_outputs[6] = packed_outputs[272:234]; correct_outputs[7] = packed_outputs[311:273]; correct_outputs[8] = packed_outputs[350:312]; correct_outputs[9] = packed_outputs[389:351]; correct_outputs[10] = packed_outputs[428:390]; correct_outputs[11] = packed_outputs[467:429]; correct_outputs[12] = packed_outputs[506:468]; correct_outputs[13] = packed_outputs[545:507]; correct_outputs[14] = packed_outputs[584:546]; correct_outputs[15] = packed_outputs[623:585]; correct_outputs[16] = packed_outputs[662:624]; correct_outputs[17] = packed_outputs[701:663]; correct_outputs[18] = packed_outputs[740:702]; correct_outputs[19] = packed_outputs[779:741]; correct_outputs[20] = packed_outputs[818:780]; correct_outputs[21] = packed_outputs[857:819]; correct_outputs[22] = packed_outputs[896:858]; correct_outputs[23] = packed_outputs[935:897]; correct_outputs[24] = packed_outputs[974:936]; correct_outputs[25] = packed_outputs[1013:975]; correct_outputs[26] = packed_outputs[1052:1014]; correct_outputs[27] = packed_outputs[1091:1053]; correct_outputs[28] = packed_outputs[1130:1092]; correct_outputs[29] = packed_outputs[1169:1131]; correct_outputs[30] = packed_outputs[1208:1170]; correct_outputs[31] = packed_outputs[1247:1209]; correct_outputs[32] = packed_outputs[1286:1248]; correct_outputs[33] = packed_outputs[1325:1287]; correct_outputs[34] = packed_outputs[1364:1326]; correct_outputs[35] = packed_outputs[1403:1365]; correct_outputs[36] = packed_outputs[1442:1404]; correct_outputs[37] = packed_outputs[1481:1443]; correct_outputs[38] = packed_outputs[1520:1482]; correct_outputs[39] = packed_outputs[1559:1521]; correct_outputs[40] = packed_outputs[1598:1560]; correct_outputs[41] = packed_outputs[1637:1599]; correct_outputs[42] = packed_outputs[1676:1638]; correct_outputs[43] = packed_outputs[1715:1677]; correct_outputs[44] = packed_outputs[1754:1716]; correct_outputs[45] = packed_outputs[1793:1755]; correct_outputs[46] = packed_outputs[1832:1794]; correct_outputs[47] = packed_outputs[1871:1833]; correct_outputs[48] = packed_outputs[1910:1872]; correct_outputs[49] = packed_outputs[1949:1911]; correct_outputs[50] = packed_outputs[1988:1950]; correct_outputs[51] = packed_outputs[2027:1989]; correct_outputs[52] = packed_outputs[2066:2028]; correct_outputs[53] = packed_outputs[2105:2067]; correct_outputs[54] = packed_outputs[2144:2106]; correct_outputs[55] = packed_outputs[2183:2145]; correct_outputs[56] = packed_outputs[2222:2184]; correct_outputs[57] = packed_outputs[2261:2223]; correct_outputs[58] = packed_outputs[2300:2262]; correct_outputs[59] = packed_outputs[2339:2301]; correct_outputs[60] = packed_outputs[2378:2340]; correct_outputs[61] = packed_outputs[2417:2379]; correct_outputs[62] = packed_outputs[2456:2418]; correct_outputs[63] = packed_outputs[2495:2457]; correct_outputs[64] = packed_outputs[2534:2496]; correct_outputs[65] = packed_outputs[2573:2535]; correct_outputs[66] = packed_outputs[2612:2574]; correct_outputs[67] = packed_outputs[2651:2613]; correct_outputs[68] = packed_outputs[2690:2652]; correct_outputs[69] = packed_outputs[2729:2691]; correct_outputs[70] = packed_outputs[2768:2730]; correct_outputs[71] = packed_outputs[2807:2769]; correct_outputs[72] = packed_outputs[2846:2808]; correct_outputs[73] = packed_outputs[2885:2847]; correct_outputs[74] = packed_outputs[2924:2886]; correct_outputs[75] = packed_outputs[2963:2925]; correct_outputs[76] = packed_outputs[3002:2964]; correct_outputs[77] = packed_outputs[3041:3003]; correct_outputs[78] = packed_outputs[3080:3042]; correct_outputs[79] = packed_outputs[3119:3081]; correct_outputs[80] = packed_outputs[3158:3120]; correct_outputs[81] = packed_outputs[3197:3159]; correct_outputs[82] = packed_outputs[3236:3198]; correct_outputs[83] = packed_outputs[3275:3237]; correct_outputs[84] = packed_outputs[3314:3276]; correct_outputs[85] = packed_outputs[3353:3315]; correct_outputs[86] = packed_outputs[3392:3354]; correct_outputs[87] = packed_outputs[3431:3393]; correct_outputs[88] = packed_outputs[3470:3432]; correct_outputs[89] = packed_outputs[3509:3471]; correct_outputs[90] = packed_outputs[3548:3510]; correct_outputs[91] = packed_outputs[3587:3549]; correct_outputs[92] = packed_outputs[3626:3588]; correct_outputs[93] = packed_outputs[3665:3627]; correct_outputs[94] = packed_outputs[3704:3666]; correct_outputs[95] = packed_outputs[3743:3705]; correct_outputs[96] = packed_outputs[3782:3744]; correct_outputs[97] = packed_outputs[3821:3783]; correct_outputs[98] = packed_outputs[3860:3822]; correct_outputs[99] = packed_outputs[3899:3861]; correct_outputs[100] = packed_outputs[3938:3900]; correct_outputs[101] = packed_outputs[3977:3939]; correct_outputs[102] = packed_outputs[4016:3978]; correct_outputs[103] = packed_outputs[4055:4017]; correct_outputs[104] = packed_outputs[4094:4056]; correct_outputs[105] = packed_outputs[4133:4095]; correct_outputs[106] = packed_outputs[4172:4134]; correct_outputs[107] = packed_outputs[4211:4173]; correct_outputs[108] = packed_outputs[4250:4212]; correct_outputs[109] = packed_outputs[4289:4251]; correct_outputs[110] = packed_outputs[4328:4290]; correct_outputs[111] = packed_outputs[4367:4329]; correct_outputs[112] = packed_outputs[4406:4368]; correct_outputs[113] = packed_outputs[4445:4407]; correct_outputs[114] = packed_outputs[4484:4446]; correct_outputs[115] = packed_outputs[4523:4485]; correct_outputs[116] = packed_outputs[4562:4524]; correct_outputs[117] = packed_outputs[4601:4563]; correct_outputs[118] = packed_outputs[4640:4602]; correct_outputs[119] = packed_outputs[4679:4641]; correct_outputs[120] = packed_outputs[4718:4680]; correct_outputs[121] = packed_outputs[4757:4719]; correct_outputs[122] = packed_outputs[4796:4758]; correct_outputs[123] = packed_outputs[4835:4797]; correct_outputs[124] = packed_outputs[4874:4836]; correct_outputs[125] = packed_outputs[4913:4875]; correct_outputs[126] = packed_outputs[4952:4914]; correct_outputs[127] = packed_outputs[4991:4953]; correct_outputs[128] = packed_outputs[5030:4992]; correct_outputs[129] = packed_outputs[5069:5031]; correct_outputs[130] = packed_outputs[5108:5070]; correct_outputs[131] = packed_outputs[5147:5109]; correct_outputs[132] = packed_outputs[5186:5148]; correct_outputs[133] = packed_outputs[5225:5187]; correct_outputs[134] = packed_outputs[5264:5226]; correct_outputs[135] = packed_outputs[5303:5265]; correct_outputs[136] = packed_outputs[5342:5304]; correct_outputs[137] = packed_outputs[5381:5343]; correct_outputs[138] = packed_outputs[5420:5382]; correct_outputs[139] = packed_outputs[5459:5421]; correct_outputs[140] = packed_outputs[5498:5460]; correct_outputs[141] = packed_outputs[5537:5499]; correct_outputs[142] = packed_outputs[5576:5538]; correct_outputs[143] = packed_outputs[5615:5577]; correct_outputs[144] = packed_outputs[5654:5616]; correct_outputs[145] = packed_outputs[5693:5655]; correct_outputs[146] = packed_outputs[5732:5694]; correct_outputs[147] = packed_outputs[5771:5733]; correct_outputs[148] = packed_outputs[5810:5772]; correct_outputs[149] = packed_outputs[5849:5811]; correct_outputs[150] = packed_outputs[5888:5850]; correct_outputs[151] = packed_outputs[5927:5889]; correct_outputs[152] = packed_outputs[5966:5928]; correct_outputs[153] = packed_outputs[6005:5967]; correct_outputs[154] = packed_outputs[6044:6006]; correct_outputs[155] = packed_outputs[6083:6045]; correct_outputs[156] = packed_outputs[6122:6084]; correct_outputs[157] = packed_outputs[6161:6123]; correct_outputs[158] = packed_outputs[6200:6162]; correct_outputs[159] = packed_outputs[6239:6201]; correct_outputs[160] = packed_outputs[6278:6240]; correct_outputs[161] = packed_outputs[6317:6279]; correct_outputs[162] = packed_outputs[6356:6318]; correct_outputs[163] = packed_outputs[6395:6357]; correct_outputs[164] = packed_outputs[6434:6396]; correct_outputs[165] = packed_outputs[6473:6435]; correct_outputs[166] = packed_outputs[6512:6474]; correct_outputs[167] = packed_outputs[6551:6513]; correct_outputs[168] = packed_outputs[6590:6552]; correct_outputs[169] = packed_outputs[6629:6591]; correct_outputs[170] = packed_outputs[6668:6630]; correct_outputs[171] = packed_outputs[6707:6669]; correct_outputs[172] = packed_outputs[6746:6708]; correct_outputs[173] = packed_outputs[6785:6747]; correct_outputs[174] = packed_outputs[6824:6786]; correct_outputs[175] = packed_outputs[6863:6825]; correct_outputs[176] = packed_outputs[6902:6864]; correct_outputs[177] = packed_outputs[6941:6903]; correct_outputs[178] = packed_outputs[6980:6942]; correct_outputs[179] = packed_outputs[7019:6981]; correct_outputs[180] = packed_outputs[7058:7020]; correct_outputs[181] = packed_outputs[7097:7059]; correct_outputs[182] = packed_outputs[7136:7098]; correct_outputs[183] = packed_outputs[7175:7137]; correct_outputs[184] = packed_outputs[7214:7176]; correct_outputs[185] = packed_outputs[7253:7215]; correct_outputs[186] = packed_outputs[7292:7254]; correct_outputs[187] = packed_outputs[7331:7293]; correct_outputs[188] = packed_outputs[7370:7332]; correct_outputs[189] = packed_outputs[7409:7371]; correct_outputs[190] = packed_outputs[7448:7410]; correct_outputs[191] = packed_outputs[7487:7449]; correct_outputs[192] = packed_outputs[7526:7488]; correct_outputs[193] = packed_outputs[7565:7527]; correct_outputs[194] = packed_outputs[7604:7566]; correct_outputs[195] = packed_outputs[7643:7605]; correct_outputs[196] = packed_outputs[7682:7644]; correct_outputs[197] = packed_outputs[7721:7683]; correct_outputs[198] = packed_outputs[7760:7722]; correct_outputs[199] = packed_outputs[7799:7761]; correct_outputs[200] = packed_outputs[7838:7800]; correct_outputs[201] = packed_outputs[7877:7839]; correct_outputs[202] = packed_outputs[7916:7878]; correct_outputs[203] = packed_outputs[7955:7917]; correct_outputs[204] = packed_outputs[7994:7956]; correct_outputs[205] = packed_outputs[8033:7995]; correct_outputs[206] = packed_outputs[8072:8034]; correct_outputs[207] = packed_outputs[8111:8073]; correct_outputs[208] = packed_outputs[8150:8112]; correct_outputs[209] = packed_outputs[8189:8151]; correct_outputs[210] = packed_outputs[8228:8190]; correct_outputs[211] = packed_outputs[8267:8229]; correct_outputs[212] = packed_outputs[8306:8268]; correct_outputs[213] = packed_outputs[8345:8307]; correct_outputs[214] = packed_outputs[8384:8346]; correct_outputs[215] = packed_outputs[8423:8385]; correct_outputs[216] = packed_outputs[8462:8424]; correct_outputs[217] = packed_outputs[8501:8463]; correct_outputs[218] = packed_outputs[8540:8502]; correct_outputs[219] = packed_outputs[8579:8541]; correct_outputs[220] = packed_outputs[8618:8580]; correct_outputs[221] = packed_outputs[8657:8619]; correct_outputs[222] = packed_outputs[8696:8658]; correct_outputs[223] = packed_outputs[8735:8697]; correct_outputs[224] = packed_outputs[8774:8736]; correct_outputs[225] = packed_outputs[8813:8775]; correct_outputs[226] = packed_outputs[8852:8814]; correct_outputs[227] = packed_outputs[8891:8853]; correct_outputs[228] = packed_outputs[8930:8892]; correct_outputs[229] = packed_outputs[8969:8931]; correct_outputs[230] = packed_outputs[9008:8970]; correct_outputs[231] = packed_outputs[9047:9009]; correct_outputs[232] = packed_outputs[9086:9048]; correct_outputs[233] = packed_outputs[9125:9087]; correct_outputs[234] = packed_outputs[9164:9126]; correct_outputs[235] = packed_outputs[9203:9165]; correct_outputs[236] = packed_outputs[9242:9204]; correct_outputs[237] = packed_outputs[9281:9243]; correct_outputs[238] = packed_outputs[9320:9282]; correct_outputs[239] = packed_outputs[9359:9321]; correct_outputs[240] = packed_outputs[9398:9360]; correct_outputs[241] = packed_outputs[9437:9399]; correct_outputs[242] = packed_outputs[9476:9438]; correct_outputs[243] = packed_outputs[9515:9477]; correct_outputs[244] = packed_outputs[9554:9516]; correct_outputs[245] = packed_outputs[9593:9555]; correct_outputs[246] = packed_outputs[9632:9594]; correct_outputs[247] = packed_outputs[9671:9633]; correct_outputs[248] = packed_outputs[9710:9672]; correct_outputs[249] = packed_outputs[9749:9711]; correct_outputs[250] = packed_outputs[9788:9750]; correct_outputs[251] = packed_outputs[9827:9789]; correct_outputs[252] = packed_outputs[9866:9828]; correct_outputs[253] = packed_outputs[9905:9867]; correct_outputs[254] = packed_outputs[9944:9906]; correct_outputs[255] = packed_outputs[9983:9945]; correct_outputs[256] = packed_outputs[10022:9984]; correct_outputs[257] = packed_outputs[10061:10023]; correct_outputs[258] = packed_outputs[10100:10062]; correct_outputs[259] = packed_outputs[10139:10101]; correct_outputs[260] = packed_outputs[10178:10140]; correct_outputs[261] = packed_outputs[10217:10179]; correct_outputs[262] = packed_outputs[10256:10218]; correct_outputs[263] = packed_outputs[10295:10257]; correct_outputs[264] = packed_outputs[10334:10296]; correct_outputs[265] = packed_outputs[10373:10335]; correct_outputs[266] = packed_outputs[10412:10374]; correct_outputs[267] = packed_outputs[10451:10413]; correct_outputs[268] = packed_outputs[10490:10452]; correct_outputs[269] = packed_outputs[10529:10491]; correct_outputs[270] = packed_outputs[10568:10530]; correct_outputs[271] = packed_outputs[10607:10569]; correct_outputs[272] = packed_outputs[10646:10608]; correct_outputs[273] = packed_outputs[10685:10647]; correct_outputs[274] = packed_outputs[10724:10686]; correct_outputs[275] = packed_outputs[10763:10725]; correct_outputs[276] = packed_outputs[10802:10764]; correct_outputs[277] = packed_outputs[10841:10803]; correct_outputs[278] = packed_outputs[10880:10842]; correct_outputs[279] = packed_outputs[10919:10881]; correct_outputs[280] = packed_outputs[10958:10920]; correct_outputs[281] = packed_outputs[10997:10959]; correct_outputs[282] = packed_outputs[11036:10998]; correct_outputs[283] = packed_outputs[11075:11037]; correct_outputs[284] = packed_outputs[11114:11076]; correct_outputs[285] = packed_outputs[11153:11115]; correct_outputs[286] = packed_outputs[11192:11154]; correct_outputs[287] = packed_outputs[11231:11193]; correct_outputs[288] = packed_outputs[11270:11232]; correct_outputs[289] = packed_outputs[11309:11271]; correct_outputs[290] = packed_outputs[11348:11310]; correct_outputs[291] = packed_outputs[11387:11349]; correct_outputs[292] = packed_outputs[11426:11388]; correct_outputs[293] = packed_outputs[11465:11427]; correct_outputs[294] = packed_outputs[11504:11466]; correct_outputs[295] = packed_outputs[11543:11505]; correct_outputs[296] = packed_outputs[11582:11544]; correct_outputs[297] = packed_outputs[11621:11583]; correct_outputs[298] = packed_outputs[11660:11622]; correct_outputs[299] = packed_outputs[11699:11661]; correct_outputs[300] = packed_outputs[11738:11700]; correct_outputs[301] = packed_outputs[11777:11739]; correct_outputs[302] = packed_outputs[11816:11778]; correct_outputs[303] = packed_outputs[11855:11817]; correct_outputs[304] = packed_outputs[11894:11856]; correct_outputs[305] = packed_outputs[11933:11895]; correct_outputs[306] = packed_outputs[11972:11934]; correct_outputs[307] = packed_outputs[12011:11973]; correct_outputs[308] = packed_outputs[12050:12012]; correct_outputs[309] = packed_outputs[12089:12051]; correct_outputs[310] = packed_outputs[12128:12090]; correct_outputs[311] = packed_outputs[12167:12129]; correct_outputs[312] = packed_outputs[12206:12168]; correct_outputs[313] = packed_outputs[12245:12207]; correct_outputs[314] = packed_outputs[12284:12246]; correct_outputs[315] = packed_outputs[12323:12285]; correct_outputs[316] = packed_outputs[12362:12324]; correct_outputs[317] = packed_outputs[12401:12363]; correct_outputs[318] = packed_outputs[12440:12402]; correct_outputs[319] = packed_outputs[12479:12441]; correct_outputs[320] = packed_outputs[12518:12480]; correct_outputs[321] = packed_outputs[12557:12519]; correct_outputs[322] = packed_outputs[12596:12558]; correct_outputs[323] = packed_outputs[12635:12597]; correct_outputs[324] = packed_outputs[12674:12636]; correct_outputs[325] = packed_outputs[12713:12675]; correct_outputs[326] = packed_outputs[12752:12714]; correct_outputs[327] = packed_outputs[12791:12753]; correct_outputs[328] = packed_outputs[12830:12792]; correct_outputs[329] = packed_outputs[12869:12831]; correct_outputs[330] = packed_outputs[12908:12870]; correct_outputs[331] = packed_outputs[12947:12909]; correct_outputs[332] = packed_outputs[12986:12948]; correct_outputs[333] = packed_outputs[13025:12987]; correct_outputs[334] = packed_outputs[13064:13026]; correct_outputs[335] = packed_outputs[13103:13065]; correct_outputs[336] = packed_outputs[13142:13104]; correct_outputs[337] = packed_outputs[13181:13143]; correct_outputs[338] = packed_outputs[13220:13182]; correct_outputs[339] = packed_outputs[13259:13221]; correct_outputs[340] = packed_outputs[13298:13260]; correct_outputs[341] = packed_outputs[13337:13299]; correct_outputs[342] = packed_outputs[13376:13338]; correct_outputs[343] = packed_outputs[13415:13377]; correct_outputs[344] = packed_outputs[13454:13416]; correct_outputs[345] = packed_outputs[13493:13455]; correct_outputs[346] = packed_outputs[13532:13494]; correct_outputs[347] = packed_outputs[13571:13533]; correct_outputs[348] = packed_outputs[13610:13572]; correct_outputs[349] = packed_outputs[13649:13611]; correct_outputs[350] = packed_outputs[13688:13650]; correct_outputs[351] = packed_outputs[13727:13689]; correct_outputs[352] = packed_outputs[13766:13728]; correct_outputs[353] = packed_outputs[13805:13767]; correct_outputs[354] = packed_outputs[13844:13806]; correct_outputs[355] = packed_outputs[13883:13845]; correct_outputs[356] = packed_outputs[13922:13884]; correct_outputs[357] = packed_outputs[13961:13923]; correct_outputs[358] = packed_outputs[14000:13962]; correct_outputs[359] = packed_outputs[14039:14001]; correct_outputs[360] = packed_outputs[14078:14040]; correct_outputs[361] = packed_outputs[14117:14079]; correct_outputs[362] = packed_outputs[14156:14118]; correct_outputs[363] = packed_outputs[14195:14157]; correct_outputs[364] = packed_outputs[14234:14196]; correct_outputs[365] = packed_outputs[14273:14235]; correct_outputs[366] = packed_outputs[14312:14274]; correct_outputs[367] = packed_outputs[14351:14313]; correct_outputs[368] = packed_outputs[14390:14352]; correct_outputs[369] = packed_outputs[14429:14391]; correct_outputs[370] = packed_outputs[14468:14430]; correct_outputs[371] = packed_outputs[14507:14469]; correct_outputs[372] = packed_outputs[14546:14508]; correct_outputs[373] = packed_outputs[14585:14547]; correct_outputs[374] = packed_outputs[14624:14586]; correct_outputs[375] = packed_outputs[14663:14625]; correct_outputs[376] = packed_outputs[14702:14664]; correct_outputs[377] = packed_outputs[14741:14703]; correct_outputs[378] = packed_outputs[14780:14742]; correct_outputs[379] = packed_outputs[14819:14781]; correct_outputs[380] = packed_outputs[14858:14820]; correct_outputs[381] = packed_outputs[14897:14859]; correct_outputs[382] = packed_outputs[14936:14898]; correct_outputs[383] = packed_outputs[14975:14937]; correct_outputs[384] = packed_outputs[15014:14976]; correct_outputs[385] = packed_outputs[15053:15015]; correct_outputs[386] = packed_outputs[15092:15054]; correct_outputs[387] = packed_outputs[15131:15093]; correct_outputs[388] = packed_outputs[15170:15132]; correct_outputs[389] = packed_outputs[15209:15171]; correct_outputs[390] = packed_outputs[15248:15210]; correct_outputs[391] = packed_outputs[15287:15249]; correct_outputs[392] = packed_outputs[15326:15288]; correct_outputs[393] = packed_outputs[15365:15327]; correct_outputs[394] = packed_outputs[15404:15366]; correct_outputs[395] = packed_outputs[15443:15405]; correct_outputs[396] = packed_outputs[15482:15444]; correct_outputs[397] = packed_outputs[15521:15483]; correct_outputs[398] = packed_outputs[15560:15522]; correct_outputs[399] = packed_outputs[15599:15561]; 
end

// END PASTE CODE

fir UUT(.clk(clk), .rst(rst), .ena(shift_ena), .sample(next_sample), .out(out));

// logic signed [38:0] diff_2;
// logic signed [38:0] diff_1;
// logic signed [38:0] diff1;
// logic signed [38:0] diff2;

always_comb begin : simulated_output
  next_sample = samples[counter];
  correct_out = correct_outputs[counter];
  diff = correct_out - out;
  // diff1 = correct_outputs[counter + 1] - out;
  // diff2 = correct_outputs[counter + 2] - out;
  // diff_1 = correct_outputs[counter - 1] - out;
  // diff_2 = correct_outputs[counter - 2] - out;
end

task print_io;
  // $display("%d %b | %b (%b), diff = %d, %d, %d, %d, %d", counter, next_sample, out, correct_out, diff, diff1, diff2, diff_1, diff_2);
  $display("%d %b | %b (%b), diff = %d", counter, next_sample, out, correct_out, diff);
endtask

integer i;
// 2) the test cases - initial blocks are like programming, not hardware
initial begin
  $dumpfile("test_fir.fst");
  $dumpvars(0, UUT);
  
  $display("Checking all inputs.");
  $display("counter, next_sample, out, correct_out");
  shift_ena = 1'b1;
  #1 clk = 1'b0;
  #1 rst = 1'b1;
  #1 clk = 1'b1;
  #1 rst = 1'b0;

  for (i = 0; i < 400; i = i + 1) begin
    #1 clk = 1'b0;
    #1 counter = i;
    #1 clk = 1'b1;
    #1 print_io();
  end

  # 1;
  if (errors !== 0) begin
    $display("---------------------------------------------------------------");
    $display("-- FAILURE                                                   --");
    $display("---------------------------------------------------------------");
    $display(" %d failures found, try again!", errors);
  end else begin
    $display("---------------------------------------------------------------");
    $display("-- SUCCESS                                                   --");
    $display("---------------------------------------------------------------");
  end
  $finish;
end

always @(counter) begin
  #1;
  assert(out === correct_out) else begin
    // $display("  ERROR: mux out should be %b, is %b", out, correct_out);
    errors = errors + 1;
  end
end

endmodule
