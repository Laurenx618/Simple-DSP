`timescale 1ns/1ps
`default_nettype none

module test_fir;
int errors = 0;

logic rst;
logic clk;
logic shift_ena;
logic [15:0] next_sample;
logic [38:0] out;

integer counter;
logic [38:0] correct_out;

// integer samples [399:0];
// time correct_outputs [399:0];

// integer test[7:0] = '{26, 40, 32, 18, 50, 0, 20, 12};

logic [6399:0] packed_samples;
always_comb packed_samples = {16'sd72200, 16'sd90564, 16'sd84560, 16'sd69249, 16'sd61880, 16'sd62782, 16'sd68570, 16'sd81332, 16'sd94609, 16'sd90928, 16'sd68018, 16'sd50830, 16'sd60149, 16'sd82167, 16'sd87989, 16'sd73243, 16'sd57675, 16'sd52510, 16'sd51258, 16'sd50538, 16'sd55715, 16'sd62361, 16'sd55290, 16'sd34526, 16'sd21916, 16'sd30203, 16'sd43308, 16'sd41391, 16'sd29511, 16'sd24186, 16'sd25102, 16'sd21159, 16'sd15385, 16'sd20309, 16'sd32017, 16'sd32431, 16'sd19016, 16'sd10144, 16'sd15839, 16'sd24055, 16'sd24052, 16'sd23069, 16'sd27703, 16'sd27689, 16'sd15133, 16'sd4539, 16'sd13068, 16'sd30953, 16'sd33500, 16'sd17189, 16'sd2083, 16'sd285, 16'sd3981, 16'sd6034, 16'sd9679, 16'sd11979, 16'sd273, -16'sd23603, -16'sd35588, -16'sd21648, -16'sd2036, -16'sd5176, -16'sd29137, -16'sd48491, -16'sd50637, -16'sd44308, -16'sd37770, -16'sd31734, -16'sd32851, -16'sd49977, -16'sd72284, -16'sd73939, -16'sd50365, -16'sd30053, -16'sd37381, -16'sd60647, -16'sd72199, -16'sd65414, -16'sd53639, -16'sd44751, -16'sd38284, -16'sd39913, -16'sd54997, -16'sd69881, -16'sd63259, -16'sd39071, -16'sd26151, -16'sd38780, -16'sd58084, -16'sd61974, -16'sd53912, -16'sd48621, -16'sd47214, -16'sd44413, -16'sd46378, -16'sd60060, -16'sd73625, -16'sd69785, -16'sd54562, -16'sd50811, -16'sd63842, -16'sd75484, -16'sd74877, -16'sd72574, -16'sd76889, -16'sd78285, -16'sd69917, -16'sd64582, -16'sd74259, -16'sd87402, -16'sd85623, -16'sd72412, -16'sd65348, -16'sd67389, -16'sd67272, -16'sd63934, -16'sd67143, -16'sd73576, -16'sd66462, -16'sd45189, -16'sd32841, -16'sd43136, -16'sd58894, -16'sd57455, -16'sd41512, -16'sd28654, -16'sd24131, -16'sd22699, -16'sd26315, -16'sd37964, -16'sd44563, -16'sd30123, -16'sd5142, 16'sd803, -16'sd19940, -16'sd41141, -16'sd39240, -16'sd21920, -16'sd9767, -16'sd8381, -16'sd12995, -16'sd23823, -16'sd38106, -16'sd39920, -16'sd19831, 16'sd2908, 16'sd475, -16'sd24053, -16'sd39415, -16'sd28863, -16'sd8252, 16'sd2297, 16'sd2573, -16'sd201, -16'sd6524, -16'sd13625, -16'sd7621, 16'sd15524, 16'sd34841, 16'sd29802, 16'sd11438, 16'sd7624, 16'sd23788, 16'sd40026, 16'sd44162, 16'sd44243, 16'sd46388, 16'sd44119, 16'sd37264, 16'sd39659, 16'sd55722, 16'sd67626, 16'sd60806, 16'sd47107, 16'sd45709, 16'sd53871, 16'sd56109, 16'sd52444, 16'sd54953, 16'sd61471, 16'sd57052, 16'sd42284, 16'sd36632, 16'sd47857, 16'sd59327, 16'sd56694, 16'sd47929, 16'sd45194, 16'sd44894, 16'sd41038, 16'sd42346, 16'sd56495, 16'sd69175, 16'sd61417, 16'sd41542, 16'sd36777, 16'sd54359, 16'sd73163, 16'sd76108, 16'sd69276, 16'sd63563, 16'sd59005, 16'sd56979, 16'sd67306, 16'sd88359, 16'sd97492, 16'sd80076, 16'sd55594, 16'sd54275, 16'sd75927, 16'sd93004, 16'sd89641, 16'sd75718, 16'sd63820, 16'sd55526, 16'sd53710, 16'sd64926, 16'sd80774, 16'sd78167, 16'sd51607, 16'sd27679, 16'sd31352, 16'sd51987, 16'sd60659, 16'sd49618, 16'sd34417, 16'sd25441, 16'sd20213, 16'sd20188, 16'sd30859, 16'sd43109, 16'sd37752, 16'sd15623, 16'sd2352, 16'sd13036, 16'sd30861, 16'sd33647, 16'sd24387, 16'sd19070, 16'sd19062, 16'sd16004, 16'sd13667, 16'sd21902, 16'sd33662, 16'sd31294, 16'sd15725, 16'sd7297, 16'sd14211, 16'sd21534, 16'sd18099, 16'sd13075, 16'sd14897, 16'sd13663, 16'sd496, -16'sd11880, -16'sd7586, 16'sd4738, 16'sd3732, -16'sd12195, -16'sd25387, -16'sd28104, -16'sd29130, -16'sd31812, -16'sd28790, -16'sd22976, -16'sd30556, -16'sd52992, -16'sd66681, -16'sd55179, -16'sd35119, -16'sd33006, -16'sd49211, -16'sd63552, -16'sd66259, -16'sd62817, -16'sd55393, -16'sd42605, -16'sd35234, -16'sd47762, -16'sd70903, -16'sd75619, -16'sd52851, -16'sd28929, -16'sd29994, -16'sd49024, -16'sd62122, -16'sd61365, -16'sd54274, -16'sd44363, -16'sd33227, -16'sd32705, -16'sd51548, -16'sd73528, -16'sd72226, -16'sd48969, -16'sd34001, -16'sd45172, -16'sd66553, -16'sd75999, -16'sd73381, -16'sd69255, -16'sd64503, -16'sd58211, -16'sd60628, -16'sd77811, -16'sd93445, -16'sd87555, -16'sd67699, -16'sd59904, -16'sd70989, -16'sd82065, -16'sd80488, -16'sd75171, -16'sd74270, -16'sd70330, -16'sd59084, -16'sd53206, -16'sd61601, -16'sd70581, -16'sd63552, -16'sd47489, -16'sd40689, -16'sd43481, -16'sd42192, -16'sd36149, -16'sd37264, -16'sd43871, -16'sd39331, -16'sd21535, -16'sd11103, -16'sd20502, -16'sd34650, -16'sd34814, -16'sd24749, -16'sd18246, -16'sd15960, -16'sd12598, -16'sd14486, -16'sd28329, -16'sd40490, -16'sd31319, -16'sd7952, 16'sd657, -16'sd15831, -16'sd35487, -16'sd36772, -16'sd24243, -16'sd12673, -16'sd5511, -16'sd2311, -16'sd9437, -16'sd25482, -16'sd30192, -16'sd9126, 16'sd19530, 16'sd24844, 16'sd5447, -16'sd9852, -16'sd2557, 16'sd16510, 16'sd30895, 16'sd38336, 16'sd39908, 16'sd31520, 16'sd18804, 16'sd21432, 16'sd45866, 16'sd68469, 16'sd64470, 16'sd42914, 16'sd32951, 16'sd43357, 16'sd57234, 16'sd62299, 16'sd62881, 16'sd61428, 16'sd52203, 16'sd39608, 16'sd40547, 16'sd57687, 16'sd69331, 16'sd59531, 16'sd42018, 16'sd38357, 16'sd46595, 16'sd50475, 16'sd48395, 16'sd50949, 16'sd56230, 16'sd51666, 16'sd39761, 16'sd38568, 16'sd52410, 16'sd63591, 16'sd60569, 16'sd54303, 16'sd56340, 16'sd59885, 16'sd56962, 16'sd57159};
logic [15:0] samples[0:399];
always_comb begin 
samples[0] = packed_samples[15:0]; samples[1] = packed_samples[31:16]; samples[2] = packed_samples[47:32]; samples[3] = packed_samples[63:48]; samples[4] = packed_samples[79:64]; samples[5] = packed_samples[95:80]; samples[6] = packed_samples[111:96]; samples[7] = packed_samples[127:112]; samples[8] = packed_samples[143:128]; samples[9] = packed_samples[159:144]; samples[10] = packed_samples[175:160]; samples[11] = packed_samples[191:176]; samples[12] = packed_samples[207:192]; samples[13] = packed_samples[223:208]; samples[14] = packed_samples[239:224]; samples[15] = packed_samples[255:240]; samples[16] = packed_samples[271:256]; samples[17] = packed_samples[287:272]; samples[18] = packed_samples[303:288]; samples[19] = packed_samples[319:304]; samples[20] = packed_samples[335:320]; samples[21] = packed_samples[351:336]; samples[22] = packed_samples[367:352]; samples[23] = packed_samples[383:368]; samples[24] = packed_samples[399:384]; samples[25] = packed_samples[415:400]; samples[26] = packed_samples[431:416]; samples[27] = packed_samples[447:432]; samples[28] = packed_samples[463:448]; samples[29] = packed_samples[479:464]; samples[30] = packed_samples[495:480]; samples[31] = packed_samples[511:496]; samples[32] = packed_samples[527:512]; samples[33] = packed_samples[543:528]; samples[34] = packed_samples[559:544]; samples[35] = packed_samples[575:560]; samples[36] = packed_samples[591:576]; samples[37] = packed_samples[607:592]; samples[38] = packed_samples[623:608]; samples[39] = packed_samples[639:624]; samples[40] = packed_samples[655:640]; samples[41] = packed_samples[671:656]; samples[42] = packed_samples[687:672]; samples[43] = packed_samples[703:688]; samples[44] = packed_samples[719:704]; samples[45] = packed_samples[735:720]; samples[46] = packed_samples[751:736]; samples[47] = packed_samples[767:752]; samples[48] = packed_samples[783:768]; samples[49] = packed_samples[799:784]; samples[50] = packed_samples[815:800]; samples[51] = packed_samples[831:816]; samples[52] = packed_samples[847:832]; samples[53] = packed_samples[863:848]; samples[54] = packed_samples[879:864]; samples[55] = packed_samples[895:880]; samples[56] = packed_samples[911:896]; samples[57] = packed_samples[927:912]; samples[58] = packed_samples[943:928]; samples[59] = packed_samples[959:944]; samples[60] = packed_samples[975:960]; samples[61] = packed_samples[991:976]; samples[62] = packed_samples[1007:992]; samples[63] = packed_samples[1023:1008]; samples[64] = packed_samples[1039:1024]; samples[65] = packed_samples[1055:1040]; samples[66] = packed_samples[1071:1056]; samples[67] = packed_samples[1087:1072]; samples[68] = packed_samples[1103:1088]; samples[69] = packed_samples[1119:1104]; samples[70] = packed_samples[1135:1120]; samples[71] = packed_samples[1151:1136]; samples[72] = packed_samples[1167:1152]; samples[73] = packed_samples[1183:1168]; samples[74] = packed_samples[1199:1184]; samples[75] = packed_samples[1215:1200]; samples[76] = packed_samples[1231:1216]; samples[77] = packed_samples[1247:1232]; samples[78] = packed_samples[1263:1248]; samples[79] = packed_samples[1279:1264]; samples[80] = packed_samples[1295:1280]; samples[81] = packed_samples[1311:1296]; samples[82] = packed_samples[1327:1312]; samples[83] = packed_samples[1343:1328]; samples[84] = packed_samples[1359:1344]; samples[85] = packed_samples[1375:1360]; samples[86] = packed_samples[1391:1376]; samples[87] = packed_samples[1407:1392]; samples[88] = packed_samples[1423:1408]; samples[89] = packed_samples[1439:1424]; samples[90] = packed_samples[1455:1440]; samples[91] = packed_samples[1471:1456]; samples[92] = packed_samples[1487:1472]; samples[93] = packed_samples[1503:1488]; samples[94] = packed_samples[1519:1504]; samples[95] = packed_samples[1535:1520]; samples[96] = packed_samples[1551:1536]; samples[97] = packed_samples[1567:1552]; samples[98] = packed_samples[1583:1568]; samples[99] = packed_samples[1599:1584]; samples[100] = packed_samples[1615:1600]; samples[101] = packed_samples[1631:1616]; samples[102] = packed_samples[1647:1632]; samples[103] = packed_samples[1663:1648]; samples[104] = packed_samples[1679:1664]; samples[105] = packed_samples[1695:1680]; samples[106] = packed_samples[1711:1696]; samples[107] = packed_samples[1727:1712]; samples[108] = packed_samples[1743:1728]; samples[109] = packed_samples[1759:1744]; samples[110] = packed_samples[1775:1760]; samples[111] = packed_samples[1791:1776]; samples[112] = packed_samples[1807:1792]; samples[113] = packed_samples[1823:1808]; samples[114] = packed_samples[1839:1824]; samples[115] = packed_samples[1855:1840]; samples[116] = packed_samples[1871:1856]; samples[117] = packed_samples[1887:1872]; samples[118] = packed_samples[1903:1888]; samples[119] = packed_samples[1919:1904]; samples[120] = packed_samples[1935:1920]; samples[121] = packed_samples[1951:1936]; samples[122] = packed_samples[1967:1952]; samples[123] = packed_samples[1983:1968]; samples[124] = packed_samples[1999:1984]; samples[125] = packed_samples[2015:2000]; samples[126] = packed_samples[2031:2016]; samples[127] = packed_samples[2047:2032]; samples[128] = packed_samples[2063:2048]; samples[129] = packed_samples[2079:2064]; samples[130] = packed_samples[2095:2080]; samples[131] = packed_samples[2111:2096]; samples[132] = packed_samples[2127:2112]; samples[133] = packed_samples[2143:2128]; samples[134] = packed_samples[2159:2144]; samples[135] = packed_samples[2175:2160]; samples[136] = packed_samples[2191:2176]; samples[137] = packed_samples[2207:2192]; samples[138] = packed_samples[2223:2208]; samples[139] = packed_samples[2239:2224]; samples[140] = packed_samples[2255:2240]; samples[141] = packed_samples[2271:2256]; samples[142] = packed_samples[2287:2272]; samples[143] = packed_samples[2303:2288]; samples[144] = packed_samples[2319:2304]; samples[145] = packed_samples[2335:2320]; samples[146] = packed_samples[2351:2336]; samples[147] = packed_samples[2367:2352]; samples[148] = packed_samples[2383:2368]; samples[149] = packed_samples[2399:2384]; samples[150] = packed_samples[2415:2400]; samples[151] = packed_samples[2431:2416]; samples[152] = packed_samples[2447:2432]; samples[153] = packed_samples[2463:2448]; samples[154] = packed_samples[2479:2464]; samples[155] = packed_samples[2495:2480]; samples[156] = packed_samples[2511:2496]; samples[157] = packed_samples[2527:2512]; samples[158] = packed_samples[2543:2528]; samples[159] = packed_samples[2559:2544]; samples[160] = packed_samples[2575:2560]; samples[161] = packed_samples[2591:2576]; samples[162] = packed_samples[2607:2592]; samples[163] = packed_samples[2623:2608]; samples[164] = packed_samples[2639:2624]; samples[165] = packed_samples[2655:2640]; samples[166] = packed_samples[2671:2656]; samples[167] = packed_samples[2687:2672]; samples[168] = packed_samples[2703:2688]; samples[169] = packed_samples[2719:2704]; samples[170] = packed_samples[2735:2720]; samples[171] = packed_samples[2751:2736]; samples[172] = packed_samples[2767:2752]; samples[173] = packed_samples[2783:2768]; samples[174] = packed_samples[2799:2784]; samples[175] = packed_samples[2815:2800]; samples[176] = packed_samples[2831:2816]; samples[177] = packed_samples[2847:2832]; samples[178] = packed_samples[2863:2848]; samples[179] = packed_samples[2879:2864]; samples[180] = packed_samples[2895:2880]; samples[181] = packed_samples[2911:2896]; samples[182] = packed_samples[2927:2912]; samples[183] = packed_samples[2943:2928]; samples[184] = packed_samples[2959:2944]; samples[185] = packed_samples[2975:2960]; samples[186] = packed_samples[2991:2976]; samples[187] = packed_samples[3007:2992]; samples[188] = packed_samples[3023:3008]; samples[189] = packed_samples[3039:3024]; samples[190] = packed_samples[3055:3040]; samples[191] = packed_samples[3071:3056]; samples[192] = packed_samples[3087:3072]; samples[193] = packed_samples[3103:3088]; samples[194] = packed_samples[3119:3104]; samples[195] = packed_samples[3135:3120]; samples[196] = packed_samples[3151:3136]; samples[197] = packed_samples[3167:3152]; samples[198] = packed_samples[3183:3168]; samples[199] = packed_samples[3199:3184]; samples[200] = packed_samples[3215:3200]; samples[201] = packed_samples[3231:3216]; samples[202] = packed_samples[3247:3232]; samples[203] = packed_samples[3263:3248]; samples[204] = packed_samples[3279:3264]; samples[205] = packed_samples[3295:3280]; samples[206] = packed_samples[3311:3296]; samples[207] = packed_samples[3327:3312]; samples[208] = packed_samples[3343:3328]; samples[209] = packed_samples[3359:3344]; samples[210] = packed_samples[3375:3360]; samples[211] = packed_samples[3391:3376]; samples[212] = packed_samples[3407:3392]; samples[213] = packed_samples[3423:3408]; samples[214] = packed_samples[3439:3424]; samples[215] = packed_samples[3455:3440]; samples[216] = packed_samples[3471:3456]; samples[217] = packed_samples[3487:3472]; samples[218] = packed_samples[3503:3488]; samples[219] = packed_samples[3519:3504]; samples[220] = packed_samples[3535:3520]; samples[221] = packed_samples[3551:3536]; samples[222] = packed_samples[3567:3552]; samples[223] = packed_samples[3583:3568]; samples[224] = packed_samples[3599:3584]; samples[225] = packed_samples[3615:3600]; samples[226] = packed_samples[3631:3616]; samples[227] = packed_samples[3647:3632]; samples[228] = packed_samples[3663:3648]; samples[229] = packed_samples[3679:3664]; samples[230] = packed_samples[3695:3680]; samples[231] = packed_samples[3711:3696]; samples[232] = packed_samples[3727:3712]; samples[233] = packed_samples[3743:3728]; samples[234] = packed_samples[3759:3744]; samples[235] = packed_samples[3775:3760]; samples[236] = packed_samples[3791:3776]; samples[237] = packed_samples[3807:3792]; samples[238] = packed_samples[3823:3808]; samples[239] = packed_samples[3839:3824]; samples[240] = packed_samples[3855:3840]; samples[241] = packed_samples[3871:3856]; samples[242] = packed_samples[3887:3872]; samples[243] = packed_samples[3903:3888]; samples[244] = packed_samples[3919:3904]; samples[245] = packed_samples[3935:3920]; samples[246] = packed_samples[3951:3936]; samples[247] = packed_samples[3967:3952]; samples[248] = packed_samples[3983:3968]; samples[249] = packed_samples[3999:3984]; samples[250] = packed_samples[4015:4000]; samples[251] = packed_samples[4031:4016]; samples[252] = packed_samples[4047:4032]; samples[253] = packed_samples[4063:4048]; samples[254] = packed_samples[4079:4064]; samples[255] = packed_samples[4095:4080]; samples[256] = packed_samples[4111:4096]; samples[257] = packed_samples[4127:4112]; samples[258] = packed_samples[4143:4128]; samples[259] = packed_samples[4159:4144]; samples[260] = packed_samples[4175:4160]; samples[261] = packed_samples[4191:4176]; samples[262] = packed_samples[4207:4192]; samples[263] = packed_samples[4223:4208]; samples[264] = packed_samples[4239:4224]; samples[265] = packed_samples[4255:4240]; samples[266] = packed_samples[4271:4256]; samples[267] = packed_samples[4287:4272]; samples[268] = packed_samples[4303:4288]; samples[269] = packed_samples[4319:4304]; samples[270] = packed_samples[4335:4320]; samples[271] = packed_samples[4351:4336]; samples[272] = packed_samples[4367:4352]; samples[273] = packed_samples[4383:4368]; samples[274] = packed_samples[4399:4384]; samples[275] = packed_samples[4415:4400]; samples[276] = packed_samples[4431:4416]; samples[277] = packed_samples[4447:4432]; samples[278] = packed_samples[4463:4448]; samples[279] = packed_samples[4479:4464]; samples[280] = packed_samples[4495:4480]; samples[281] = packed_samples[4511:4496]; samples[282] = packed_samples[4527:4512]; samples[283] = packed_samples[4543:4528]; samples[284] = packed_samples[4559:4544]; samples[285] = packed_samples[4575:4560]; samples[286] = packed_samples[4591:4576]; samples[287] = packed_samples[4607:4592]; samples[288] = packed_samples[4623:4608]; samples[289] = packed_samples[4639:4624]; samples[290] = packed_samples[4655:4640]; samples[291] = packed_samples[4671:4656]; samples[292] = packed_samples[4687:4672]; samples[293] = packed_samples[4703:4688]; samples[294] = packed_samples[4719:4704]; samples[295] = packed_samples[4735:4720]; samples[296] = packed_samples[4751:4736]; samples[297] = packed_samples[4767:4752]; samples[298] = packed_samples[4783:4768]; samples[299] = packed_samples[4799:4784]; samples[300] = packed_samples[4815:4800]; samples[301] = packed_samples[4831:4816]; samples[302] = packed_samples[4847:4832]; samples[303] = packed_samples[4863:4848]; samples[304] = packed_samples[4879:4864]; samples[305] = packed_samples[4895:4880]; samples[306] = packed_samples[4911:4896]; samples[307] = packed_samples[4927:4912]; samples[308] = packed_samples[4943:4928]; samples[309] = packed_samples[4959:4944]; samples[310] = packed_samples[4975:4960]; samples[311] = packed_samples[4991:4976]; samples[312] = packed_samples[5007:4992]; samples[313] = packed_samples[5023:5008]; samples[314] = packed_samples[5039:5024]; samples[315] = packed_samples[5055:5040]; samples[316] = packed_samples[5071:5056]; samples[317] = packed_samples[5087:5072]; samples[318] = packed_samples[5103:5088]; samples[319] = packed_samples[5119:5104]; samples[320] = packed_samples[5135:5120]; samples[321] = packed_samples[5151:5136]; samples[322] = packed_samples[5167:5152]; samples[323] = packed_samples[5183:5168]; samples[324] = packed_samples[5199:5184]; samples[325] = packed_samples[5215:5200]; samples[326] = packed_samples[5231:5216]; samples[327] = packed_samples[5247:5232]; samples[328] = packed_samples[5263:5248]; samples[329] = packed_samples[5279:5264]; samples[330] = packed_samples[5295:5280]; samples[331] = packed_samples[5311:5296]; samples[332] = packed_samples[5327:5312]; samples[333] = packed_samples[5343:5328]; samples[334] = packed_samples[5359:5344]; samples[335] = packed_samples[5375:5360]; samples[336] = packed_samples[5391:5376]; samples[337] = packed_samples[5407:5392]; samples[338] = packed_samples[5423:5408]; samples[339] = packed_samples[5439:5424]; samples[340] = packed_samples[5455:5440]; samples[341] = packed_samples[5471:5456]; samples[342] = packed_samples[5487:5472]; samples[343] = packed_samples[5503:5488]; samples[344] = packed_samples[5519:5504]; samples[345] = packed_samples[5535:5520]; samples[346] = packed_samples[5551:5536]; samples[347] = packed_samples[5567:5552]; samples[348] = packed_samples[5583:5568]; samples[349] = packed_samples[5599:5584]; samples[350] = packed_samples[5615:5600]; samples[351] = packed_samples[5631:5616]; samples[352] = packed_samples[5647:5632]; samples[353] = packed_samples[5663:5648]; samples[354] = packed_samples[5679:5664]; samples[355] = packed_samples[5695:5680]; samples[356] = packed_samples[5711:5696]; samples[357] = packed_samples[5727:5712]; samples[358] = packed_samples[5743:5728]; samples[359] = packed_samples[5759:5744]; samples[360] = packed_samples[5775:5760]; samples[361] = packed_samples[5791:5776]; samples[362] = packed_samples[5807:5792]; samples[363] = packed_samples[5823:5808]; samples[364] = packed_samples[5839:5824]; samples[365] = packed_samples[5855:5840]; samples[366] = packed_samples[5871:5856]; samples[367] = packed_samples[5887:5872]; samples[368] = packed_samples[5903:5888]; samples[369] = packed_samples[5919:5904]; samples[370] = packed_samples[5935:5920]; samples[371] = packed_samples[5951:5936]; samples[372] = packed_samples[5967:5952]; samples[373] = packed_samples[5983:5968]; samples[374] = packed_samples[5999:5984]; samples[375] = packed_samples[6015:6000]; samples[376] = packed_samples[6031:6016]; samples[377] = packed_samples[6047:6032]; samples[378] = packed_samples[6063:6048]; samples[379] = packed_samples[6079:6064]; samples[380] = packed_samples[6095:6080]; samples[381] = packed_samples[6111:6096]; samples[382] = packed_samples[6127:6112]; samples[383] = packed_samples[6143:6128]; samples[384] = packed_samples[6159:6144]; samples[385] = packed_samples[6175:6160]; samples[386] = packed_samples[6191:6176]; samples[387] = packed_samples[6207:6192]; samples[388] = packed_samples[6223:6208]; samples[389] = packed_samples[6239:6224]; samples[390] = packed_samples[6255:6240]; samples[391] = packed_samples[6271:6256]; samples[392] = packed_samples[6287:6272]; samples[393] = packed_samples[6303:6288]; samples[394] = packed_samples[6319:6304]; samples[395] = packed_samples[6335:6320]; samples[396] = packed_samples[6351:6336]; samples[397] = packed_samples[6367:6352]; samples[398] = packed_samples[6383:6368]; samples[399] = packed_samples[6399:6384]; 
end

logic [15599:0] packed_outputs;
always_comb packed_outputs = {-39'sd680344, -39'sd1249027, -39'sd729189, 39'sd1604747, 39'sd5510102, 39'sd9517597, 39'sd11225695, 39'sd8257649, -39'sd193474, -39'sd12036352, -39'sd22348746, -39'sd25225238, -39'sd16561402, 39'sd3491148, 39'sd29339678, 39'sd50756621, 39'sd56169119, 39'sd37863337, -39'sd3036453, -39'sd54530355, -39'sd96273242, -39'sd106458679, -39'sd71194131, 39'sd6905391, 39'sd105038314, 39'sd184675544, 39'sd204221742, 39'sd136129330, -39'sd17532302, -39'sd217019524, -39'sd388544939, -39'sd440467321, -39'sd288384022, 39'sd118584483, 39'sd779191628, 39'sd1635563348, 39'sd2584669271, 39'sd3502834615, 39'sd4276283405, 39'sd4828391583, 39'sd5135234107, 39'sd5225309636, 39'sd5164910509, 39'sd5034855787, 39'sd4906215322, 39'sd4822415457, 39'sd4792702820, 39'sd4797583806, 39'sd4802346973, 39'sd4772542544, 39'sd4686012972, 39'sd4538371451, 39'sd4341351108, 39'sd4115844880, 39'sd3883239565, 39'sd3658740346, 39'sd3448620675, 39'sd3251205834, 39'sd3060318524, 39'sd2869667374, 39'sd2676482228, 39'sd2482894746, 39'sd2294752510, 39'sd2119050508, 39'sd1961578198, 39'sd1825613808, 39'sd1711726412, 39'sd1618520094, 39'sd1543913620, 39'sd1486144420, 39'sd1443869537, 39'sd1415644487, 39'sd1399583439, 39'sd1393463392, 39'sd1395334482, 39'sd1401729440, 39'sd1409349257, 39'sd1415045527, 39'sd1415850343, 39'sd1408712506, 39'sd1390536666, 39'sd1358577801, 39'sd1310619698, 39'sd1244769489, 39'sd1159378250, 39'sd1053322259, 39'sd926173231, 39'sd777959263, 39'sd608969735, 39'sd420003136, 39'sd212650657, -39'sd10913061, -39'sd248349975, -39'sd497174709, -39'sd754468102, -39'sd1016886292, -39'sd1281003119, -39'sd1543457205, -39'sd1800804872, -39'sd2049565754, -39'sd2286582415, -39'sd2509171523, -39'sd2714850626, -39'sd2901186975, -39'sd3066152536, -39'sd3208510380, -39'sd3327686683, -39'sd3423422757, -39'sd3495798444, -39'sd3545508820, -39'sd3573857267, -39'sd3582500163, -39'sd3573432974, -39'sd3549199200, -39'sd3512799363, -39'sd3467265063, -39'sd3415496545, -39'sd3360558259, -39'sd3305839757, -39'sd3254699227, -39'sd3210064736, -39'sd3174496235, -39'sd3150405255, -39'sd3139924554, -39'sd3144621437, -39'sd3165540193, -39'sd3203424056, -39'sd3258607773, -39'sd3330685529, -39'sd3418535575, -39'sd3520714474, -39'sd3635599843, -39'sd3761099757, -39'sd3894502523, -39'sd4032789086, -39'sd4172935175, -39'sd4311800463, -39'sd4445976249, -39'sd4572031477, -39'sd4686852519, -39'sd4787584312, -39'sd4871399638, -39'sd4935642688, -39'sd4978220836, -39'sd4997660593, -39'sd4992829193, -39'sd4962900316, -39'sd4907672195, -39'sd4827680589, -39'sd4723895831, -39'sd4597532075, -39'sd4450290469, -39'sd4284564647, -39'sd4103175270, -39'sd3909004474, -39'sd3705042483, -39'sd3494606792, -39'sd3281207797, -39'sd3068202212, -39'sd2858757240, -39'sd2656048658, -39'sd2463150213, -39'sd2282625860, -39'sd2116424109, -39'sd1966200130, -39'sd1833456980, -39'sd1719204103, -39'sd1623656724, -39'sd1546414429, -39'sd1486748438, -39'sd1443526511, -39'sd1415026426, -39'sd1399085387, -39'sd1393370079, -39'sd1395295928, -39'sd1401790068, -39'sd1409464270, -39'sd1415100177, -39'sd1415786123, -39'sd1408603216, -39'sd1390497512, -39'sd1358629108, -39'sd1310688480, -39'sd1244798133, -39'sd1159370150, -39'sd1053293395, -39'sd926128433, -39'sd777925344, -39'sd608988455, -39'sd420066199, -39'sd212691504, 39'sd10934638, 39'sd248397668, 39'sd497197646, 39'sd754467482, 39'sd1016883018, 39'sd1280984437, 39'sd1543410748, 39'sd1800774184, 39'sd2049604907, 39'sd2286664496, 39'sd2509206000, 39'sd2714798709, 39'sd2901106593, 39'sd3066118168, 39'sd3208537826, 39'sd3327749115, 39'sd3423485907, 39'sd3495816523, 39'sd3545443790, 39'sd3573745968, 39'sd3582455603, 39'sd3573520576, 39'sd3549337687, 39'sd3512842807, 39'sd3467172225, 39'sd3415367382, 39'sd3360510300, 39'sd3305899952, 39'sd3254812416, 39'sd3210148441, 39'sd3174480190, 39'sd3150283010, 39'sd3139794481, 39'sd3144618918, 39'sd3165684339, 39'sd3203571636, 39'sd3258606538, 39'sd3330545359, 39'sd3418403248, 39'sd3520704793, 39'sd3635700554, 39'sd3761219909, 39'sd3894553703, 39'sd4032729101, 39'sd4172800524, 39'sd4311707126, 39'sd4446025029, 39'sd4572184634, 39'sd4686953560, 39'sd4787531885, 39'sd4871260505, 39'sd4935560374, 39'sd4978254569, 39'sd4997755454, 39'sd4992904798, 39'sd4962912248, 39'sd4907612851, 39'sd4827586364, 39'sd4723847872, 39'sd4597586417, 39'sd4450397588, 39'sd4284611380, 39'sd4103119995, 39'sd3908921125, 39'sd3705015107, 39'sd3494635095, 39'sd3281244745, 39'sd3068229565, 39'sd2858776599, 39'sd2656040446, 39'sd2463101764, 39'sd2282578193, 39'sd2116432099, 39'sd1966254228, 39'sd1833495929, 39'sd1719199916, 39'sd1623634864, 39'sd1546392840, 39'sd1486718012, 39'sd1443502820, 39'sd1415054996, 39'sd1399162709, 39'sd1393414651, 39'sd1395245950, 39'sd1401693470, 39'sd1409422554, 39'sd1415147310, 39'sd1415868176, 39'sd1408654856, 39'sd1390489290, 39'sd1358560455, 39'sd1310596159, 39'sd1244764317, 39'sd1159451978, 39'sd1053428891, 39'sd926175129, 39'sd777824466, 39'sd608843488, 39'sd420023277, 39'sd212780111, -39'sd10808148, -39'sd248337736, -39'sd497242634, -39'sd754585812, -39'sd1016987672, -39'sd1280976052, -39'sd1543274751, -39'sd1800632613, -39'sd2049607436, -39'sd2286814417, -39'sd2509347418, -39'sd2714794080, -39'sd2900978726, -39'sd3065996868, -39'sd3208517740, -39'sd3327830782, -39'sd3423605111, -39'sd3495883247, -39'sd3545392107, -39'sd3573606695, -39'sd3582359936, -39'sd3573571599, -39'sd3549483501, -39'sd3512929988, -39'sd3467123377, -39'sd3415252806, -39'sd3360442234, -39'sd3305916345, -39'sd3254880663, -39'sd3210220934, -39'sd3174510140, -39'sd3150237439, -39'sd3139701628, -39'sd3144568920, -39'sd3165732296, -39'sd3203662281, -39'sd3258641808, -39'sd3330505867, -39'sd3418351351, -39'sd3520685062, -39'sd3635700760, -39'sd3761228064, -39'sd3894584255, -39'sd4032772495, -39'sd4172807431, -39'sd4311658050, -39'sd4445970880, -39'sd4572181051, -39'sd4686991143, -39'sd4787567414, -39'sd4871279918, -39'sd4935566636, -39'sd4978229092, -39'sd4997691858, -39'sd4992859933, -39'sd4962953888, -39'sd4907714681, -39'sd4827638970, -39'sd4723791830, -39'sd4597483119, -39'sd4450347189, -39'sd4284646649, -39'sd4103203019, -39'sd3908994940, -39'sd3705026191, -39'sd3494555712, -39'sd3281124440, -39'sd3068186830, -39'sd2858875461, -39'sd2656191254, -39'sd2463146118, -39'sd2282471426, -39'sd2116288505, -39'sd1966208814, -39'sd1833573049, -39'sd1719323701, -39'sd1623710967, -39'sd1546362187, -39'sd1486591395, -39'sd1443380596, -39'sd1415061729, -39'sd1399309517, -39'sd1393558099, -39'sd1395236836, -39'sd1401547290, -39'sd1409293513, -39'sd1415149926, -39'sd1415976828, -39'sd1408766703, -39'sd1390523934, -39'sd1358496187, -39'sd1310475479, -39'sd1244686307, -39'sd1159499955, -39'sd1053567883, -39'sd926264615, -39'sd777772732, -39'sd608714815, -39'sd419953035, -39'sd212818149, 39'sd10723054, 39'sd248279976, 39'sd497238088, 39'sd754630761, 39'sd1017059437, 39'sd1281019096, 39'sd1543239093, 39'sd1800546637, 39'sd2049562238};
logic [38:0] correct_outputs[0:399];
always_comb begin
correct_outputs[0] = packed_outputs[38:0]; correct_outputs[1] = packed_outputs[77:39]; correct_outputs[2] = packed_outputs[116:78]; correct_outputs[3] = packed_outputs[155:117]; correct_outputs[4] = packed_outputs[194:156]; correct_outputs[5] = packed_outputs[233:195]; correct_outputs[6] = packed_outputs[272:234]; correct_outputs[7] = packed_outputs[311:273]; correct_outputs[8] = packed_outputs[350:312]; correct_outputs[9] = packed_outputs[389:351]; correct_outputs[10] = packed_outputs[428:390]; correct_outputs[11] = packed_outputs[467:429]; correct_outputs[12] = packed_outputs[506:468]; correct_outputs[13] = packed_outputs[545:507]; correct_outputs[14] = packed_outputs[584:546]; correct_outputs[15] = packed_outputs[623:585]; correct_outputs[16] = packed_outputs[662:624]; correct_outputs[17] = packed_outputs[701:663]; correct_outputs[18] = packed_outputs[740:702]; correct_outputs[19] = packed_outputs[779:741]; correct_outputs[20] = packed_outputs[818:780]; correct_outputs[21] = packed_outputs[857:819]; correct_outputs[22] = packed_outputs[896:858]; correct_outputs[23] = packed_outputs[935:897]; correct_outputs[24] = packed_outputs[974:936]; correct_outputs[25] = packed_outputs[1013:975]; correct_outputs[26] = packed_outputs[1052:1014]; correct_outputs[27] = packed_outputs[1091:1053]; correct_outputs[28] = packed_outputs[1130:1092]; correct_outputs[29] = packed_outputs[1169:1131]; correct_outputs[30] = packed_outputs[1208:1170]; correct_outputs[31] = packed_outputs[1247:1209]; correct_outputs[32] = packed_outputs[1286:1248]; correct_outputs[33] = packed_outputs[1325:1287]; correct_outputs[34] = packed_outputs[1364:1326]; correct_outputs[35] = packed_outputs[1403:1365]; correct_outputs[36] = packed_outputs[1442:1404]; correct_outputs[37] = packed_outputs[1481:1443]; correct_outputs[38] = packed_outputs[1520:1482]; correct_outputs[39] = packed_outputs[1559:1521]; correct_outputs[40] = packed_outputs[1598:1560]; correct_outputs[41] = packed_outputs[1637:1599]; correct_outputs[42] = packed_outputs[1676:1638]; correct_outputs[43] = packed_outputs[1715:1677]; correct_outputs[44] = packed_outputs[1754:1716]; correct_outputs[45] = packed_outputs[1793:1755]; correct_outputs[46] = packed_outputs[1832:1794]; correct_outputs[47] = packed_outputs[1871:1833]; correct_outputs[48] = packed_outputs[1910:1872]; correct_outputs[49] = packed_outputs[1949:1911]; correct_outputs[50] = packed_outputs[1988:1950]; correct_outputs[51] = packed_outputs[2027:1989]; correct_outputs[52] = packed_outputs[2066:2028]; correct_outputs[53] = packed_outputs[2105:2067]; correct_outputs[54] = packed_outputs[2144:2106]; correct_outputs[55] = packed_outputs[2183:2145]; correct_outputs[56] = packed_outputs[2222:2184]; correct_outputs[57] = packed_outputs[2261:2223]; correct_outputs[58] = packed_outputs[2300:2262]; correct_outputs[59] = packed_outputs[2339:2301]; correct_outputs[60] = packed_outputs[2378:2340]; correct_outputs[61] = packed_outputs[2417:2379]; correct_outputs[62] = packed_outputs[2456:2418]; correct_outputs[63] = packed_outputs[2495:2457]; correct_outputs[64] = packed_outputs[2534:2496]; correct_outputs[65] = packed_outputs[2573:2535]; correct_outputs[66] = packed_outputs[2612:2574]; correct_outputs[67] = packed_outputs[2651:2613]; correct_outputs[68] = packed_outputs[2690:2652]; correct_outputs[69] = packed_outputs[2729:2691]; correct_outputs[70] = packed_outputs[2768:2730]; correct_outputs[71] = packed_outputs[2807:2769]; correct_outputs[72] = packed_outputs[2846:2808]; correct_outputs[73] = packed_outputs[2885:2847]; correct_outputs[74] = packed_outputs[2924:2886]; correct_outputs[75] = packed_outputs[2963:2925]; correct_outputs[76] = packed_outputs[3002:2964]; correct_outputs[77] = packed_outputs[3041:3003]; correct_outputs[78] = packed_outputs[3080:3042]; correct_outputs[79] = packed_outputs[3119:3081]; correct_outputs[80] = packed_outputs[3158:3120]; correct_outputs[81] = packed_outputs[3197:3159]; correct_outputs[82] = packed_outputs[3236:3198]; correct_outputs[83] = packed_outputs[3275:3237]; correct_outputs[84] = packed_outputs[3314:3276]; correct_outputs[85] = packed_outputs[3353:3315]; correct_outputs[86] = packed_outputs[3392:3354]; correct_outputs[87] = packed_outputs[3431:3393]; correct_outputs[88] = packed_outputs[3470:3432]; correct_outputs[89] = packed_outputs[3509:3471]; correct_outputs[90] = packed_outputs[3548:3510]; correct_outputs[91] = packed_outputs[3587:3549]; correct_outputs[92] = packed_outputs[3626:3588]; correct_outputs[93] = packed_outputs[3665:3627]; correct_outputs[94] = packed_outputs[3704:3666]; correct_outputs[95] = packed_outputs[3743:3705]; correct_outputs[96] = packed_outputs[3782:3744]; correct_outputs[97] = packed_outputs[3821:3783]; correct_outputs[98] = packed_outputs[3860:3822]; correct_outputs[99] = packed_outputs[3899:3861]; correct_outputs[100] = packed_outputs[3938:3900]; correct_outputs[101] = packed_outputs[3977:3939]; correct_outputs[102] = packed_outputs[4016:3978]; correct_outputs[103] = packed_outputs[4055:4017]; correct_outputs[104] = packed_outputs[4094:4056]; correct_outputs[105] = packed_outputs[4133:4095]; correct_outputs[106] = packed_outputs[4172:4134]; correct_outputs[107] = packed_outputs[4211:4173]; correct_outputs[108] = packed_outputs[4250:4212]; correct_outputs[109] = packed_outputs[4289:4251]; correct_outputs[110] = packed_outputs[4328:4290]; correct_outputs[111] = packed_outputs[4367:4329]; correct_outputs[112] = packed_outputs[4406:4368]; correct_outputs[113] = packed_outputs[4445:4407]; correct_outputs[114] = packed_outputs[4484:4446]; correct_outputs[115] = packed_outputs[4523:4485]; correct_outputs[116] = packed_outputs[4562:4524]; correct_outputs[117] = packed_outputs[4601:4563]; correct_outputs[118] = packed_outputs[4640:4602]; correct_outputs[119] = packed_outputs[4679:4641]; correct_outputs[120] = packed_outputs[4718:4680]; correct_outputs[121] = packed_outputs[4757:4719]; correct_outputs[122] = packed_outputs[4796:4758]; correct_outputs[123] = packed_outputs[4835:4797]; correct_outputs[124] = packed_outputs[4874:4836]; correct_outputs[125] = packed_outputs[4913:4875]; correct_outputs[126] = packed_outputs[4952:4914]; correct_outputs[127] = packed_outputs[4991:4953]; correct_outputs[128] = packed_outputs[5030:4992]; correct_outputs[129] = packed_outputs[5069:5031]; correct_outputs[130] = packed_outputs[5108:5070]; correct_outputs[131] = packed_outputs[5147:5109]; correct_outputs[132] = packed_outputs[5186:5148]; correct_outputs[133] = packed_outputs[5225:5187]; correct_outputs[134] = packed_outputs[5264:5226]; correct_outputs[135] = packed_outputs[5303:5265]; correct_outputs[136] = packed_outputs[5342:5304]; correct_outputs[137] = packed_outputs[5381:5343]; correct_outputs[138] = packed_outputs[5420:5382]; correct_outputs[139] = packed_outputs[5459:5421]; correct_outputs[140] = packed_outputs[5498:5460]; correct_outputs[141] = packed_outputs[5537:5499]; correct_outputs[142] = packed_outputs[5576:5538]; correct_outputs[143] = packed_outputs[5615:5577]; correct_outputs[144] = packed_outputs[5654:5616]; correct_outputs[145] = packed_outputs[5693:5655]; correct_outputs[146] = packed_outputs[5732:5694]; correct_outputs[147] = packed_outputs[5771:5733]; correct_outputs[148] = packed_outputs[5810:5772]; correct_outputs[149] = packed_outputs[5849:5811]; correct_outputs[150] = packed_outputs[5888:5850]; correct_outputs[151] = packed_outputs[5927:5889]; correct_outputs[152] = packed_outputs[5966:5928]; correct_outputs[153] = packed_outputs[6005:5967]; correct_outputs[154] = packed_outputs[6044:6006]; correct_outputs[155] = packed_outputs[6083:6045]; correct_outputs[156] = packed_outputs[6122:6084]; correct_outputs[157] = packed_outputs[6161:6123]; correct_outputs[158] = packed_outputs[6200:6162]; correct_outputs[159] = packed_outputs[6239:6201]; correct_outputs[160] = packed_outputs[6278:6240]; correct_outputs[161] = packed_outputs[6317:6279]; correct_outputs[162] = packed_outputs[6356:6318]; correct_outputs[163] = packed_outputs[6395:6357]; correct_outputs[164] = packed_outputs[6434:6396]; correct_outputs[165] = packed_outputs[6473:6435]; correct_outputs[166] = packed_outputs[6512:6474]; correct_outputs[167] = packed_outputs[6551:6513]; correct_outputs[168] = packed_outputs[6590:6552]; correct_outputs[169] = packed_outputs[6629:6591]; correct_outputs[170] = packed_outputs[6668:6630]; correct_outputs[171] = packed_outputs[6707:6669]; correct_outputs[172] = packed_outputs[6746:6708]; correct_outputs[173] = packed_outputs[6785:6747]; correct_outputs[174] = packed_outputs[6824:6786]; correct_outputs[175] = packed_outputs[6863:6825]; correct_outputs[176] = packed_outputs[6902:6864]; correct_outputs[177] = packed_outputs[6941:6903]; correct_outputs[178] = packed_outputs[6980:6942]; correct_outputs[179] = packed_outputs[7019:6981]; correct_outputs[180] = packed_outputs[7058:7020]; correct_outputs[181] = packed_outputs[7097:7059]; correct_outputs[182] = packed_outputs[7136:7098]; correct_outputs[183] = packed_outputs[7175:7137]; correct_outputs[184] = packed_outputs[7214:7176]; correct_outputs[185] = packed_outputs[7253:7215]; correct_outputs[186] = packed_outputs[7292:7254]; correct_outputs[187] = packed_outputs[7331:7293]; correct_outputs[188] = packed_outputs[7370:7332]; correct_outputs[189] = packed_outputs[7409:7371]; correct_outputs[190] = packed_outputs[7448:7410]; correct_outputs[191] = packed_outputs[7487:7449]; correct_outputs[192] = packed_outputs[7526:7488]; correct_outputs[193] = packed_outputs[7565:7527]; correct_outputs[194] = packed_outputs[7604:7566]; correct_outputs[195] = packed_outputs[7643:7605]; correct_outputs[196] = packed_outputs[7682:7644]; correct_outputs[197] = packed_outputs[7721:7683]; correct_outputs[198] = packed_outputs[7760:7722]; correct_outputs[199] = packed_outputs[7799:7761]; correct_outputs[200] = packed_outputs[7838:7800]; correct_outputs[201] = packed_outputs[7877:7839]; correct_outputs[202] = packed_outputs[7916:7878]; correct_outputs[203] = packed_outputs[7955:7917]; correct_outputs[204] = packed_outputs[7994:7956]; correct_outputs[205] = packed_outputs[8033:7995]; correct_outputs[206] = packed_outputs[8072:8034]; correct_outputs[207] = packed_outputs[8111:8073]; correct_outputs[208] = packed_outputs[8150:8112]; correct_outputs[209] = packed_outputs[8189:8151]; correct_outputs[210] = packed_outputs[8228:8190]; correct_outputs[211] = packed_outputs[8267:8229]; correct_outputs[212] = packed_outputs[8306:8268]; correct_outputs[213] = packed_outputs[8345:8307]; correct_outputs[214] = packed_outputs[8384:8346]; correct_outputs[215] = packed_outputs[8423:8385]; correct_outputs[216] = packed_outputs[8462:8424]; correct_outputs[217] = packed_outputs[8501:8463]; correct_outputs[218] = packed_outputs[8540:8502]; correct_outputs[219] = packed_outputs[8579:8541]; correct_outputs[220] = packed_outputs[8618:8580]; correct_outputs[221] = packed_outputs[8657:8619]; correct_outputs[222] = packed_outputs[8696:8658]; correct_outputs[223] = packed_outputs[8735:8697]; correct_outputs[224] = packed_outputs[8774:8736]; correct_outputs[225] = packed_outputs[8813:8775]; correct_outputs[226] = packed_outputs[8852:8814]; correct_outputs[227] = packed_outputs[8891:8853]; correct_outputs[228] = packed_outputs[8930:8892]; correct_outputs[229] = packed_outputs[8969:8931]; correct_outputs[230] = packed_outputs[9008:8970]; correct_outputs[231] = packed_outputs[9047:9009]; correct_outputs[232] = packed_outputs[9086:9048]; correct_outputs[233] = packed_outputs[9125:9087]; correct_outputs[234] = packed_outputs[9164:9126]; correct_outputs[235] = packed_outputs[9203:9165]; correct_outputs[236] = packed_outputs[9242:9204]; correct_outputs[237] = packed_outputs[9281:9243]; correct_outputs[238] = packed_outputs[9320:9282]; correct_outputs[239] = packed_outputs[9359:9321]; correct_outputs[240] = packed_outputs[9398:9360]; correct_outputs[241] = packed_outputs[9437:9399]; correct_outputs[242] = packed_outputs[9476:9438]; correct_outputs[243] = packed_outputs[9515:9477]; correct_outputs[244] = packed_outputs[9554:9516]; correct_outputs[245] = packed_outputs[9593:9555]; correct_outputs[246] = packed_outputs[9632:9594]; correct_outputs[247] = packed_outputs[9671:9633]; correct_outputs[248] = packed_outputs[9710:9672]; correct_outputs[249] = packed_outputs[9749:9711]; correct_outputs[250] = packed_outputs[9788:9750]; correct_outputs[251] = packed_outputs[9827:9789]; correct_outputs[252] = packed_outputs[9866:9828]; correct_outputs[253] = packed_outputs[9905:9867]; correct_outputs[254] = packed_outputs[9944:9906]; correct_outputs[255] = packed_outputs[9983:9945]; correct_outputs[256] = packed_outputs[10022:9984]; correct_outputs[257] = packed_outputs[10061:10023]; correct_outputs[258] = packed_outputs[10100:10062]; correct_outputs[259] = packed_outputs[10139:10101]; correct_outputs[260] = packed_outputs[10178:10140]; correct_outputs[261] = packed_outputs[10217:10179]; correct_outputs[262] = packed_outputs[10256:10218]; correct_outputs[263] = packed_outputs[10295:10257]; correct_outputs[264] = packed_outputs[10334:10296]; correct_outputs[265] = packed_outputs[10373:10335]; correct_outputs[266] = packed_outputs[10412:10374]; correct_outputs[267] = packed_outputs[10451:10413]; correct_outputs[268] = packed_outputs[10490:10452]; correct_outputs[269] = packed_outputs[10529:10491]; correct_outputs[270] = packed_outputs[10568:10530]; correct_outputs[271] = packed_outputs[10607:10569]; correct_outputs[272] = packed_outputs[10646:10608]; correct_outputs[273] = packed_outputs[10685:10647]; correct_outputs[274] = packed_outputs[10724:10686]; correct_outputs[275] = packed_outputs[10763:10725]; correct_outputs[276] = packed_outputs[10802:10764]; correct_outputs[277] = packed_outputs[10841:10803]; correct_outputs[278] = packed_outputs[10880:10842]; correct_outputs[279] = packed_outputs[10919:10881]; correct_outputs[280] = packed_outputs[10958:10920]; correct_outputs[281] = packed_outputs[10997:10959]; correct_outputs[282] = packed_outputs[11036:10998]; correct_outputs[283] = packed_outputs[11075:11037]; correct_outputs[284] = packed_outputs[11114:11076]; correct_outputs[285] = packed_outputs[11153:11115]; correct_outputs[286] = packed_outputs[11192:11154]; correct_outputs[287] = packed_outputs[11231:11193]; correct_outputs[288] = packed_outputs[11270:11232]; correct_outputs[289] = packed_outputs[11309:11271]; correct_outputs[290] = packed_outputs[11348:11310]; correct_outputs[291] = packed_outputs[11387:11349]; correct_outputs[292] = packed_outputs[11426:11388]; correct_outputs[293] = packed_outputs[11465:11427]; correct_outputs[294] = packed_outputs[11504:11466]; correct_outputs[295] = packed_outputs[11543:11505]; correct_outputs[296] = packed_outputs[11582:11544]; correct_outputs[297] = packed_outputs[11621:11583]; correct_outputs[298] = packed_outputs[11660:11622]; correct_outputs[299] = packed_outputs[11699:11661]; correct_outputs[300] = packed_outputs[11738:11700]; correct_outputs[301] = packed_outputs[11777:11739]; correct_outputs[302] = packed_outputs[11816:11778]; correct_outputs[303] = packed_outputs[11855:11817]; correct_outputs[304] = packed_outputs[11894:11856]; correct_outputs[305] = packed_outputs[11933:11895]; correct_outputs[306] = packed_outputs[11972:11934]; correct_outputs[307] = packed_outputs[12011:11973]; correct_outputs[308] = packed_outputs[12050:12012]; correct_outputs[309] = packed_outputs[12089:12051]; correct_outputs[310] = packed_outputs[12128:12090]; correct_outputs[311] = packed_outputs[12167:12129]; correct_outputs[312] = packed_outputs[12206:12168]; correct_outputs[313] = packed_outputs[12245:12207]; correct_outputs[314] = packed_outputs[12284:12246]; correct_outputs[315] = packed_outputs[12323:12285]; correct_outputs[316] = packed_outputs[12362:12324]; correct_outputs[317] = packed_outputs[12401:12363]; correct_outputs[318] = packed_outputs[12440:12402]; correct_outputs[319] = packed_outputs[12479:12441]; correct_outputs[320] = packed_outputs[12518:12480]; correct_outputs[321] = packed_outputs[12557:12519]; correct_outputs[322] = packed_outputs[12596:12558]; correct_outputs[323] = packed_outputs[12635:12597]; correct_outputs[324] = packed_outputs[12674:12636]; correct_outputs[325] = packed_outputs[12713:12675]; correct_outputs[326] = packed_outputs[12752:12714]; correct_outputs[327] = packed_outputs[12791:12753]; correct_outputs[328] = packed_outputs[12830:12792]; correct_outputs[329] = packed_outputs[12869:12831]; correct_outputs[330] = packed_outputs[12908:12870]; correct_outputs[331] = packed_outputs[12947:12909]; correct_outputs[332] = packed_outputs[12986:12948]; correct_outputs[333] = packed_outputs[13025:12987]; correct_outputs[334] = packed_outputs[13064:13026]; correct_outputs[335] = packed_outputs[13103:13065]; correct_outputs[336] = packed_outputs[13142:13104]; correct_outputs[337] = packed_outputs[13181:13143]; correct_outputs[338] = packed_outputs[13220:13182]; correct_outputs[339] = packed_outputs[13259:13221]; correct_outputs[340] = packed_outputs[13298:13260]; correct_outputs[341] = packed_outputs[13337:13299]; correct_outputs[342] = packed_outputs[13376:13338]; correct_outputs[343] = packed_outputs[13415:13377]; correct_outputs[344] = packed_outputs[13454:13416]; correct_outputs[345] = packed_outputs[13493:13455]; correct_outputs[346] = packed_outputs[13532:13494]; correct_outputs[347] = packed_outputs[13571:13533]; correct_outputs[348] = packed_outputs[13610:13572]; correct_outputs[349] = packed_outputs[13649:13611]; correct_outputs[350] = packed_outputs[13688:13650]; correct_outputs[351] = packed_outputs[13727:13689]; correct_outputs[352] = packed_outputs[13766:13728]; correct_outputs[353] = packed_outputs[13805:13767]; correct_outputs[354] = packed_outputs[13844:13806]; correct_outputs[355] = packed_outputs[13883:13845]; correct_outputs[356] = packed_outputs[13922:13884]; correct_outputs[357] = packed_outputs[13961:13923]; correct_outputs[358] = packed_outputs[14000:13962]; correct_outputs[359] = packed_outputs[14039:14001]; correct_outputs[360] = packed_outputs[14078:14040]; correct_outputs[361] = packed_outputs[14117:14079]; correct_outputs[362] = packed_outputs[14156:14118]; correct_outputs[363] = packed_outputs[14195:14157]; correct_outputs[364] = packed_outputs[14234:14196]; correct_outputs[365] = packed_outputs[14273:14235]; correct_outputs[366] = packed_outputs[14312:14274]; correct_outputs[367] = packed_outputs[14351:14313]; correct_outputs[368] = packed_outputs[14390:14352]; correct_outputs[369] = packed_outputs[14429:14391]; correct_outputs[370] = packed_outputs[14468:14430]; correct_outputs[371] = packed_outputs[14507:14469]; correct_outputs[372] = packed_outputs[14546:14508]; correct_outputs[373] = packed_outputs[14585:14547]; correct_outputs[374] = packed_outputs[14624:14586]; correct_outputs[375] = packed_outputs[14663:14625]; correct_outputs[376] = packed_outputs[14702:14664]; correct_outputs[377] = packed_outputs[14741:14703]; correct_outputs[378] = packed_outputs[14780:14742]; correct_outputs[379] = packed_outputs[14819:14781]; correct_outputs[380] = packed_outputs[14858:14820]; correct_outputs[381] = packed_outputs[14897:14859]; correct_outputs[382] = packed_outputs[14936:14898]; correct_outputs[383] = packed_outputs[14975:14937]; correct_outputs[384] = packed_outputs[15014:14976]; correct_outputs[385] = packed_outputs[15053:15015]; correct_outputs[386] = packed_outputs[15092:15054]; correct_outputs[387] = packed_outputs[15131:15093]; correct_outputs[388] = packed_outputs[15170:15132]; correct_outputs[389] = packed_outputs[15209:15171]; correct_outputs[390] = packed_outputs[15248:15210]; correct_outputs[391] = packed_outputs[15287:15249]; correct_outputs[392] = packed_outputs[15326:15288]; correct_outputs[393] = packed_outputs[15365:15327]; correct_outputs[394] = packed_outputs[15404:15366]; correct_outputs[395] = packed_outputs[15443:15405]; correct_outputs[396] = packed_outputs[15482:15444]; correct_outputs[397] = packed_outputs[15521:15483]; correct_outputs[398] = packed_outputs[15560:15522]; correct_outputs[399] = packed_outputs[15599:15561]; 
end


// // integer xyzzy[7:0] = '{26, 40, 32, 18, 50, 0, 20, 12};

// logic [15:0] samples [399:0] = '{72200, 90564, 84560, 69249, 61880, 62782, 68570, 81332, 94609, 90928, 68018, 50830, 60149, 82167, 87989, 73243, 57675, 52510, 51258, 50538, 55715, 62361, 55290, 34526, 21916, 30203, 43308, 41391, 29511, 24186, 25102, 21159, 15385, 20309, 32017, 32431, 19016, 10144, 15839, 24055, 24052, 23069, 27703, 27689, 15133, 4539, 13068, 30953, 33500, 17189, 2083, 285, 3981, 6034, 9679, 11979, 273, -23603, -35588, -21648, -2036, -5176, -29137, -48491, -50637, -44308, -37770, -31734, -32851, -49977, -72284, -73939, -50365, -30053, -37381, -60647, -72199, -65414, -53639, -44751, -38284, -39913, -54997, -69881, -63259, -39071, -26151, -38780, -58084, -61974, -53912, -48621, -47214, -44413, -46378, -60060, -73625, -69785, -54562, -50811, -63842, -75484, -74877, -72574, -76889, -78285, -69917, -64582, -74259, -87402, -85623, -72412, -65348, -67389, -67272, -63934, -67143, -73576, -66462, -45189, -32841, -43136, -58894, -57455, -41512, -28654, -24131, -22699, -26315, -37964, -44563, -30123, -5142, 803, -19940, -41141, -39240, -21920, -9767, -8381, -12995, -23823, -38106, -39920, -19831, 2908, 475, -24053, -39415, -28863, -8252, 2297, 2573, -201, -6524, -13625, -7621, 15524, 34841, 29802, 11438, 7624, 23788, 40026, 44162, 44243, 46388, 44119, 37264, 39659, 55722, 67626, 60806, 47107, 45709, 53871, 56109, 52444, 54953, 61471, 57052, 42284, 36632, 47857, 59327, 56694, 47929, 45194, 44894, 41038, 42346, 56495, 69175, 61417, 41542, 36777, 54359, 73163, 76108, 69276, 63563, 59005, 56979, 67306, 88359, 97492, 80076, 55594, 54275, 75927, 93004, 89641, 75718, 63820, 55526, 53710, 64926, 80774, 78167, 51607, 27679, 31352, 51987, 60659, 49618, 34417, 25441, 20213, 20188, 30859, 43109, 37752, 15623, 2352, 13036, 30861, 33647, 24387, 19070, 19062, 16004, 13667, 21902, 33662, 31294, 15725, 7297, 14211, 21534, 18099, 13075, 14897, 13663, 496, -11880, -7586, 4738, 3732, -12195, -25387, -28104, -29130, -31812, -28790, -22976, -30556, -52992, -66681, -55179, -35119, -33006, -49211, -63552, -66259, -62817, -55393, -42605, -35234, -47762, -70903, -75619, -52851, -28929, -29994, -49024, -62122, -61365, -54274, -44363, -33227, -32705, -51548, -73528, -72226, -48969, -34001, -45172, -66553, -75999, -73381, -69255, -64503, -58211, -60628, -77811, -93445, -87555, -67699, -59904, -70989, -82065, -80488, -75171, -74270, -70330, -59084, -53206, -61601, -70581, -63552, -47489, -40689, -43481, -42192, -36149, -37264, -43871, -39331, -21535, -11103, -20502, -34650, -34814, -24749, -18246, -15960, -12598, -14486, -28329, -40490, -31319, -7952, 657, -15831, -35487, -36772, -24243, -12673, -5511, -2311, -9437, -25482, -30192, -9126, 19530, 24844, 5447, -9852, -2557, 16510, 30895, 38336, 39908, 31520, 18804, 21432, 45866, 68469, 64470, 42914, 32951, 43357, 57234, 62299, 62881, 61428, 52203, 39608, 40547, 57687, 69331, 59531, 42018, 38357, 46595, 50475, 48395, 50949, 56230, 51666, 39761, 38568, 52410, 63591, 60569, 54303, 56340, 59885, 56962, 57159};
// logic [38:0] correct_outputs [399:0] = '{-680344, -1249027, -729189, 1604747, 5510102, 9517597, 11225695, 8257649, -193474, -12036352, -22348746, -25225238, -16561402, 3491148, 29339678, 50756621, 56169119, 37863337, -3036453, -54530355, -96273242, -106458679, -71194131, 6905391, 105038314, 184675544, 204221742, 136129330, -17532302, -217019524, -388544939, -440467321, -288384022, 118584483, 779191628, 1635563348, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2119050508, 1961578198, 1825613808, 1711726412, 1618520094, 1543913620, 1486144420, 1443869537, 1415644487, 1399583439, 1393463392, 1395334482, 1401729440, 1409349257, 1415045527, 1415850343, 1408712506, 1390536666, 1358577801, 1310619698, 1244769489, 1159378250, 1053322259, 926173231, 777959263, 608969735, 420003136, 212650657, -10913061, -248349975, -497174709, -754468102, -1016886292, -1281003119, -1543457205, -1800804872, -2049565754, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116424109, -1966200130, -1833456980, -1719204103, -1623656724, -1546414429, -1486748438, -1443526511, -1415026426, -1399085387, -1393370079, -1395295928, -1401790068, -1409464270, -1415100177, -1415786123, -1408603216, -1390497512, -1358629108, -1310688480, -1244798133, -1159370150, -1053293395, -926128433, -777925344, -608988455, -420066199, -212691504, 10934638, 248397668, 497197646, 754467482, 1016883018, 1280984437, 1543410748, 1800774184, 2049604907, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2116432099, 1966254228, 1833495929, 1719199916, 1623634864, 1546392840, 1486718012, 1443502820, 1415054996, 1399162709, 1393414651, 1395245950, 1401693470, 1409422554, 1415147310, 1415868176, 1408654856, 1390489290, 1358560455, 1310596159, 1244764317, 1159451978, 1053428891, 926175129, 777824466, 608843488, 420023277, 212780111, -10808148, -248337736, -497242634, -754585812, -1016987672, -1280976052, -1543274751, -1800632613, -2049607436, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116288505, -1966208814, -1833573049, -1719323701, -1623710967, -1546362187, -1486591395, -1443380596, -1415061729, -1399309517, -1393558099, -1395236836, -1401547290, -1409293513, -1415149926, -1415976828, -1408766703, -1390523934, -1358496187, -1310475479, -1244686307, -1159499955, -1053567883, -926264615, -777772732, -608714815, -419953035, -212818149, 10723054, 248279976, 497238088, 754630761, 1017059437, 1281019096, 1543239093, 1800546637, 2049562238};
// // always_comb samples = '{72200, 90564, 84560, 69249, 61880, 62782, 68570, 81332, 94609, 90928, 68018, 50830, 60149, 82167, 87989, 73243, 57675, 52510, 51258, 50538, 55715, 62361, 55290, 34526, 21916, 30203, 43308, 41391, 29511, 24186, 25102, 21159, 15385, 20309, 32017, 32431, 19016, 10144, 15839, 24055, 24052, 23069, 27703, 27689, 15133, 4539, 13068, 30953, 33500, 17189, 2083, 285, 3981, 6034, 9679, 11979, 273, -23603, -35588, -21648, -2036, -5176, -29137, -48491, -50637, -44308, -37770, -31734, -32851, -49977, -72284, -73939, -50365, -30053, -37381, -60647, -72199, -65414, -53639, -44751, -38284, -39913, -54997, -69881, -63259, -39071, -26151, -38780, -58084, -61974, -53912, -48621, -47214, -44413, -46378, -60060, -73625, -69785, -54562, -50811, -63842, -75484, -74877, -72574, -76889, -78285, -69917, -64582, -74259, -87402, -85623, -72412, -65348, -67389, -67272, -63934, -67143, -73576, -66462, -45189, -32841, -43136, -58894, -57455, -41512, -28654, -24131, -22699, -26315, -37964, -44563, -30123, -5142, 803, -19940, -41141, -39240, -21920, -9767, -8381, -12995, -23823, -38106, -39920, -19831, 2908, 475, -24053, -39415, -28863, -8252, 2297, 2573, -201, -6524, -13625, -7621, 15524, 34841, 29802, 11438, 7624, 23788, 40026, 44162, 44243, 46388, 44119, 37264, 39659, 55722, 67626, 60806, 47107, 45709, 53871, 56109, 52444, 54953, 61471, 57052, 42284, 36632, 47857, 59327, 56694, 47929, 45194, 44894, 41038, 42346, 56495, 69175, 61417, 41542, 36777, 54359, 73163, 76108, 69276, 63563, 59005, 56979, 67306, 88359, 97492, 80076, 55594, 54275, 75927, 93004, 89641, 75718, 63820, 55526, 53710, 64926, 80774, 78167, 51607, 27679, 31352, 51987, 60659, 49618, 34417, 25441, 20213, 20188, 30859, 43109, 37752, 15623, 2352, 13036, 30861, 33647, 24387, 19070, 19062, 16004, 13667, 21902, 33662, 31294, 15725, 7297, 14211, 21534, 18099, 13075, 14897, 13663, 496, -11880, -7586, 4738, 3732, -12195, -25387, -28104, -29130, -31812, -28790, -22976, -30556, -52992, -66681, -55179, -35119, -33006, -49211, -63552, -66259, -62817, -55393, -42605, -35234, -47762, -70903, -75619, -52851, -28929, -29994, -49024, -62122, -61365, -54274, -44363, -33227, -32705, -51548, -73528, -72226, -48969, -34001, -45172, -66553, -75999, -73381, -69255, -64503, -58211, -60628, -77811, -93445, -87555, -67699, -59904, -70989, -82065, -80488, -75171, -74270, -70330, -59084, -53206, -61601, -70581, -63552, -47489, -40689, -43481, -42192, -36149, -37264, -43871, -39331, -21535, -11103, -20502, -34650, -34814, -24749, -18246, -15960, -12598, -14486, -28329, -40490, -31319, -7952, 657, -15831, -35487, -36772, -24243, -12673, -5511, -2311, -9437, -25482, -30192, -9126, 19530, 24844, 5447, -9852, -2557, 16510, 30895, 38336, 39908, 31520, 18804, 21432, 45866, 68469, 64470, 42914, 32951, 43357, 57234, 62299, 62881, 61428, 52203, 39608, 40547, 57687, 69331, 59531, 42018, 38357, 46595, 50475, 48395, 50949, 56230, 51666, 39761, 38568, 52410, 63591, 60569, 54303, 56340, 59885, 56962, 57159};
// // always_comb correct_outputs = '{-680344, -1249027, -729189, 1604747, 5510102, 9517597, 11225695, 8257649, -193474, -12036352, -22348746, -25225238, -16561402, 3491148, 29339678, 50756621, 56169119, 37863337, -3036453, -54530355, -96273242, -106458679, -71194131, 6905391, 105038314, 184675544, 204221742, 136129330, -17532302, -217019524, -388544939, -440467321, -288384022, 118584483, 779191628, 1635563348, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2119050508, 1961578198, 1825613808, 1711726412, 1618520094, 1543913620, 1486144420, 1443869537, 1415644487, 1399583439, 1393463392, 1395334482, 1401729440, 1409349257, 1415045527, 1415850343, 1408712506, 1390536666, 1358577801, 1310619698, 1244769489, 1159378250, 1053322259, 926173231, 777959263, 608969735, 420003136, 212650657, -10913061, -248349975, -497174709, -754468102, -1016886292, -1281003119, -1543457205, -1800804872, -2049565754, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116424109, -1966200130, -1833456980, -1719204103, -1623656724, -1546414429, -1486748438, -1443526511, -1415026426, -1399085387, -1393370079, -1395295928, -1401790068, -1409464270, -1415100177, -1415786123, -1408603216, -1390497512, -1358629108, -1310688480, -1244798133, -1159370150, -1053293395, -926128433, -777925344, -608988455, -420066199, -212691504, 10934638, 248397668, 497197646, 754467482, 1016883018, 1280984437, 1543410748, 1800774184, 2049604907, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, 2116432099, 1966254228, 1833495929, 1719199916, 1623634864, 1546392840, 1486718012, 1443502820, 1415054996, 1399162709, 1393414651, 1395245950, 1401693470, 1409422554, 1415147310, 1415868176, 1408654856, 1390489290, 1358560455, 1310596159, 1244764317, 1159451978, 1053428891, 926175129, 777824466, 608843488, 420023277, 212780111, -10808148, -248337736, -497242634, -754585812, -1016987672, -1280976052, -1543274751, -1800632613, -2049607436, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2147483648, -2116288505, -1966208814, -1833573049, -1719323701, -1623710967, -1546362187, -1486591395, -1443380596, -1415061729, -1399309517, -1393558099, -1395236836, -1401547290, -1409293513, -1415149926, -1415976828, -1408766703, -1390523934, -1358496187, -1310475479, -1244686307, -1159499955, -1053567883, -926264615, -777772732, -608714815, -419953035, -212818149, 10723054, 248279976, 497238088, 754630761, 1017059437, 1281019096, 1543239093, 1800546637, 2049562238};

// module fir #(clk, rst, ena, sample, out);
fir UUT(.clk(clk), .rst(rst), .ena(shift_ena), .sample(next_sample), .out(out));

always_comb begin : simulated_output
  next_sample = samples[counter];
  correct_out = correct_outputs[counter];
end

task print_io;
  $display("%d %b | %b (%b)", counter, next_sample, out, correct_out);
endtask

integer i;
// 2) the test cases - initial blocks are like programming, not hardware
initial begin
  $dumpfile("test_fir.fst");
  $dumpvars(0, UUT);
  
  $display("Checking all inputs.");
  $display("counter, next_sample, out, correct_out");
  shift_ena = 1'b0;
  rst = 1'b1;
  #1 rst = 1'b0;
  for (i = 0; i < 400; i = i + 1) begin
    #1 clk = 1'b0;
    #1 counter = i;
    #1 clk = 1'b1;
    #1 print_io();
  end

  # 1;
  if (errors !== 0) begin
    $display("---------------------------------------------------------------");
    $display("-- FAILURE                                                   --");
    $display("---------------------------------------------------------------");
    $display(" %d failures found, try again!", errors);
  end else begin
    $display("---------------------------------------------------------------");
    $display("-- SUCCESS                                                   --");
    $display("---------------------------------------------------------------");
  end
  $finish;
end

always @(counter) begin
  #1;
  assert(out === correct_out) else begin
    // $display("  ERROR: mux out should be %b, is %b", out, correct_out);
    errors = errors + 1;
  end
end

endmodule
